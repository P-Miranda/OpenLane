`timescale 1ns / 1ps
`include "global_defines.vh"
`include "system.vh"
`include "axi.vh"
`include "xversat.vh"
`include "xdefs.vh"

module M #(
      parameter ADDR_W = `ADDR_W,
      parameter DATA_W = `DATA_W,
      parameter AXI_ADDR_W = 32
   )
   (

   input run,
   
   input [DATA_W-1:0]              in0,
   output [DATA_W-1:0]             out0,
   input [31:0]     M_Stage_sigma_constant_00_00,
   input [31:0]     M_Stage_sigma_constant_01_01,
   input [31:0]     M_Stage_sigma_constant_02_02,
   input [31:0]     M_Stage_sigma_constant_00_03,
   input [31:0]     M_Stage_sigma_constant_01_04,
   input [31:0]     M_Stage_sigma_constant_02_05,
   input [5:0]     M_buffer0_amount,
   input [5:0]     M_buffer1_amount,
   input [5:0]     M_buffer2_amount,
   input [5:0]     M_buffer3_amount,
   input [5:0]     M_buffer4_amount,
   input [5:0]     M_buffer5_amount,
   input [5:0]     M_buffer6_amount,
   input [5:0]     M_buffer7_amount,
   input [5:0]     M_buffer8_amount,
   input [5:0]     M_buffer9_amount,
   input [5:0]     M_buffer10_amount,
   input [5:0]     M_buffer11_amount,
   input [5:0]     M_buffer12_amount,
   input [5:0]     M_buffer13_amount,
   input [5:0]     M_buffer14_amount,
   input [5:0]     M_buffer15_amount,
   input [5:0]     M_buffer16_amount,
   input [5:0]     M_buffer17_amount,
   input [5:0]     M_buffer18_amount,
   input [5:0]     M_buffer19_amount,
   input [5:0]     M_buffer20_amount,
   input [5:0]     M_buffer21_amount,
   input [5:0]     M_buffer22_amount,
   input [5:0]     M_buffer23_amount,
   input [5:0]     M_buffer24_amount,
   input [5:0]     M_buffer25_amount,
   input [5:0]     M_buffer26_amount,
   input [5:0]     M_buffer27_amount,
   input [5:0]     M_buffer28_amount,
   input [5:0]     M_buffer29_amount,
   input [5:0]     M_buffer30_amount,
   input [5:0]     M_buffer31_amount,
   input [5:0]     M_buffer32_amount,
   input [5:0]     M_buffer33_amount,
   input [5:0]     M_buffer34_amount,
   input [5:0]     M_buffer35_amount,
   input [5:0]     M_buffer36_amount,
   input [5:0]     M_buffer37_amount,
   input [5:0]     M_buffer38_amount,
   input [5:0]     M_buffer39_amount,
   input [5:0]     M_buffer40_amount,
   input [5:0]     M_buffer41_amount,
   input [5:0]     M_buffer42_amount,
   input [5:0]     M_buffer43_amount,
   input [5:0]     M_buffer44_amount,
   input [5:0]     M_buffer45_amount,
   input [5:0]     M_buffer46_amount,
   input [5:0]     M_buffer47_amount,
   input [5:0]     M_buffer48_amount,
   input [5:0]     M_buffer49_amount,
   input [5:0]     M_buffer50_amount,
   input [5:0]     M_buffer51_amount,
   input [5:0]     M_buffer52_amount,
   input [5:0]     M_buffer53_amount,
   input [5:0]     M_buffer54_amount,
   input [5:0]     M_buffer55_amount,
   input [5:0]     M_buffer56_amount,
   input [5:0]     M_buffer57_amount,
   input [5:0]     M_buffer58_amount,
   input [5:0]     M_buffer59_amount,
   input [5:0]     M_buffer60_amount,
   input [5:0]     M_buffer61_amount,
   input  [31:0]                   delay0,
   input                           clk,
   input                           rst
   );

wire wor_ready;

wire [31:0] unitRdataFinal;
reg [31:0] stateRead;

wire [31:0] output_0_0 , output_1_0 , output_2_0 , output_3_0 , output_4_0 , output_5_0 , output_6_0 , output_7_0 , output_8_0 , output_9_0 , output_10_0 , output_11_0 , output_12_0 , output_13_0 , output_14_0 , output_15_0 , output_16_0 , output_17_0 , output_19_0 , output_20_0 , output_21_0 , output_22_0 , output_23_0 , output_24_0 , output_25_0 , output_26_0 , output_27_0 , output_28_0 , output_29_0 , output_30_0 , output_31_0 , output_32_0 , output_33_0 , output_34_0 , output_35_0 , output_36_0 , output_37_0 , output_38_0 , output_39_0 , output_40_0 , output_41_0 , output_42_0 , output_43_0 , output_44_0 , output_45_0 , output_46_0 , output_47_0 , output_48_0 , output_49_0 , output_50_0 , output_51_0 , output_52_0 , output_53_0 , output_54_0 , output_55_0 , output_56_0 , output_57_0 , output_58_0 , output_59_0 , output_60_0 , output_61_0 , output_62_0 , output_63_0 , output_64_0 , output_65_0 , output_66_0 , output_67_0 , output_68_0 , output_69_0 , output_70_0 , output_71_0 , output_72_0 , output_73_0 , output_74_0 , output_75_0 , output_76_0 , output_77_0 , output_78_0 , output_79_0 , output_80_0 ;

M_Stage  m0_0 (
         .out0(output_1_0),
         .in1(in0), // w
         .in0(output_43_0),
         .in2(output_44_0),
         .in3(output_45_0),
         .M_Stage_sigma_constant_00_00(M_Stage_sigma_constant_00_00),
         .M_Stage_sigma_constant_01_01(M_Stage_sigma_constant_01_01),
         .M_Stage_sigma_constant_02_02(M_Stage_sigma_constant_02_02),
         .M_Stage_sigma_constant_00_03(M_Stage_sigma_constant_00_03),
         .M_Stage_sigma_constant_01_04(M_Stage_sigma_constant_01_04),
         .M_Stage_sigma_constant_02_05(M_Stage_sigma_constant_02_05),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         M_Stage  m1_1 (
         .out0(output_2_0),
         .in1(in0), // w
         .in0(output_46_0),
         .in2(output_47_0),
         .in3(output_48_0),
         .M_Stage_sigma_constant_00_00(M_Stage_sigma_constant_00_00),
         .M_Stage_sigma_constant_01_01(M_Stage_sigma_constant_01_01),
         .M_Stage_sigma_constant_02_02(M_Stage_sigma_constant_02_02),
         .M_Stage_sigma_constant_00_03(M_Stage_sigma_constant_00_03),
         .M_Stage_sigma_constant_01_04(M_Stage_sigma_constant_01_04),
         .M_Stage_sigma_constant_02_05(M_Stage_sigma_constant_02_05),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         M_Stage  m2_2 (
         .out0(output_3_0),
         .in1(output_40_0),
         .in0(output_49_0),
         .in2(output_50_0),
         .in3(output_51_0),
         .M_Stage_sigma_constant_00_00(M_Stage_sigma_constant_00_00),
         .M_Stage_sigma_constant_01_01(M_Stage_sigma_constant_01_01),
         .M_Stage_sigma_constant_02_02(M_Stage_sigma_constant_02_02),
         .M_Stage_sigma_constant_00_03(M_Stage_sigma_constant_00_03),
         .M_Stage_sigma_constant_01_04(M_Stage_sigma_constant_01_04),
         .M_Stage_sigma_constant_02_05(M_Stage_sigma_constant_02_05),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         M_Stage  m3_3 (
         .out0(output_4_0),
         .in1(output_38_0),
         .in0(output_52_0),
         .in2(output_53_0),
         .in3(output_54_0),
         .M_Stage_sigma_constant_00_00(M_Stage_sigma_constant_00_00),
         .M_Stage_sigma_constant_01_01(M_Stage_sigma_constant_01_01),
         .M_Stage_sigma_constant_02_02(M_Stage_sigma_constant_02_02),
         .M_Stage_sigma_constant_00_03(M_Stage_sigma_constant_00_03),
         .M_Stage_sigma_constant_01_04(M_Stage_sigma_constant_01_04),
         .M_Stage_sigma_constant_02_05(M_Stage_sigma_constant_02_05),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         M_Stage  m4_4 (
         .out0(output_5_0),
         .in1(output_36_0),
         .in0(output_55_0),
         .in2(output_56_0),
         .in3(output_57_0),
         .M_Stage_sigma_constant_00_00(M_Stage_sigma_constant_00_00),
         .M_Stage_sigma_constant_01_01(M_Stage_sigma_constant_01_01),
         .M_Stage_sigma_constant_02_02(M_Stage_sigma_constant_02_02),
         .M_Stage_sigma_constant_00_03(M_Stage_sigma_constant_00_03),
         .M_Stage_sigma_constant_01_04(M_Stage_sigma_constant_01_04),
         .M_Stage_sigma_constant_02_05(M_Stage_sigma_constant_02_05),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         M_Stage  m5_5 (
         .out0(output_6_0),
         .in1(output_34_0),
         .in0(output_58_0),
         .in2(output_59_0),
         .in3(output_60_0),
         .M_Stage_sigma_constant_00_00(M_Stage_sigma_constant_00_00),
         .M_Stage_sigma_constant_01_01(M_Stage_sigma_constant_01_01),
         .M_Stage_sigma_constant_02_02(M_Stage_sigma_constant_02_02),
         .M_Stage_sigma_constant_00_03(M_Stage_sigma_constant_00_03),
         .M_Stage_sigma_constant_01_04(M_Stage_sigma_constant_01_04),
         .M_Stage_sigma_constant_02_05(M_Stage_sigma_constant_02_05),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         M_Stage  m6_6 (
         .out0(output_7_0),
         .in1(output_32_0),
         .in0(output_61_0),
         .in2(output_62_0),
         .in3(output_63_0),
         .M_Stage_sigma_constant_00_00(M_Stage_sigma_constant_00_00),
         .M_Stage_sigma_constant_01_01(M_Stage_sigma_constant_01_01),
         .M_Stage_sigma_constant_02_02(M_Stage_sigma_constant_02_02),
         .M_Stage_sigma_constant_00_03(M_Stage_sigma_constant_00_03),
         .M_Stage_sigma_constant_01_04(M_Stage_sigma_constant_01_04),
         .M_Stage_sigma_constant_02_05(M_Stage_sigma_constant_02_05),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         M_Stage  m7_7 (
         .out0(output_8_0),
         .in1(output_30_0),
         .in2(output_41_0),
         .in0(output_64_0),
         .in3(output_65_0),
         .M_Stage_sigma_constant_00_00(M_Stage_sigma_constant_00_00),
         .M_Stage_sigma_constant_01_01(M_Stage_sigma_constant_01_01),
         .M_Stage_sigma_constant_02_02(M_Stage_sigma_constant_02_02),
         .M_Stage_sigma_constant_00_03(M_Stage_sigma_constant_00_03),
         .M_Stage_sigma_constant_01_04(M_Stage_sigma_constant_01_04),
         .M_Stage_sigma_constant_02_05(M_Stage_sigma_constant_02_05),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         M_Stage  m8_8 (
         .out0(output_9_0),
         .in1(output_28_0),
         .in2(output_39_0),
         .in0(output_66_0),
         .in3(output_67_0),
         .M_Stage_sigma_constant_00_00(M_Stage_sigma_constant_00_00),
         .M_Stage_sigma_constant_01_01(M_Stage_sigma_constant_01_01),
         .M_Stage_sigma_constant_02_02(M_Stage_sigma_constant_02_02),
         .M_Stage_sigma_constant_00_03(M_Stage_sigma_constant_00_03),
         .M_Stage_sigma_constant_01_04(M_Stage_sigma_constant_01_04),
         .M_Stage_sigma_constant_02_05(M_Stage_sigma_constant_02_05),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         M_Stage  m9_9 (
         .out0(output_10_0),
         .in1(output_26_0),
         .in2(output_37_0),
         .in0(output_68_0),
         .in3(output_69_0),
         .M_Stage_sigma_constant_00_00(M_Stage_sigma_constant_00_00),
         .M_Stage_sigma_constant_01_01(M_Stage_sigma_constant_01_01),
         .M_Stage_sigma_constant_02_02(M_Stage_sigma_constant_02_02),
         .M_Stage_sigma_constant_00_03(M_Stage_sigma_constant_00_03),
         .M_Stage_sigma_constant_01_04(M_Stage_sigma_constant_01_04),
         .M_Stage_sigma_constant_02_05(M_Stage_sigma_constant_02_05),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         M_Stage  ma_10 (
         .out0(output_11_0),
         .in1(output_24_0),
         .in2(output_35_0),
         .in0(output_70_0),
         .in3(output_71_0),
         .M_Stage_sigma_constant_00_00(M_Stage_sigma_constant_00_00),
         .M_Stage_sigma_constant_01_01(M_Stage_sigma_constant_01_01),
         .M_Stage_sigma_constant_02_02(M_Stage_sigma_constant_02_02),
         .M_Stage_sigma_constant_00_03(M_Stage_sigma_constant_00_03),
         .M_Stage_sigma_constant_01_04(M_Stage_sigma_constant_01_04),
         .M_Stage_sigma_constant_02_05(M_Stage_sigma_constant_02_05),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         M_Stage  mb_11 (
         .out0(output_12_0),
         .in1(output_23_0),
         .in2(output_33_0),
         .in0(output_72_0),
         .in3(output_73_0),
         .M_Stage_sigma_constant_00_00(M_Stage_sigma_constant_00_00),
         .M_Stage_sigma_constant_01_01(M_Stage_sigma_constant_01_01),
         .M_Stage_sigma_constant_02_02(M_Stage_sigma_constant_02_02),
         .M_Stage_sigma_constant_00_03(M_Stage_sigma_constant_00_03),
         .M_Stage_sigma_constant_01_04(M_Stage_sigma_constant_01_04),
         .M_Stage_sigma_constant_02_05(M_Stage_sigma_constant_02_05),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         M_Stage  mc_12 (
         .out0(output_13_0),
         .in1(output_22_0),
         .in2(output_31_0),
         .in0(output_74_0),
         .in3(output_75_0),
         .M_Stage_sigma_constant_00_00(M_Stage_sigma_constant_00_00),
         .M_Stage_sigma_constant_01_01(M_Stage_sigma_constant_01_01),
         .M_Stage_sigma_constant_02_02(M_Stage_sigma_constant_02_02),
         .M_Stage_sigma_constant_00_03(M_Stage_sigma_constant_00_03),
         .M_Stage_sigma_constant_01_04(M_Stage_sigma_constant_01_04),
         .M_Stage_sigma_constant_02_05(M_Stage_sigma_constant_02_05),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         M_Stage  md_13 (
         .out0(output_14_0),
         .in1(output_21_0),
         .in2(output_29_0),
         .in0(output_76_0),
         .in3(output_77_0),
         .M_Stage_sigma_constant_00_00(M_Stage_sigma_constant_00_00),
         .M_Stage_sigma_constant_01_01(M_Stage_sigma_constant_01_01),
         .M_Stage_sigma_constant_02_02(M_Stage_sigma_constant_02_02),
         .M_Stage_sigma_constant_00_03(M_Stage_sigma_constant_00_03),
         .M_Stage_sigma_constant_01_04(M_Stage_sigma_constant_01_04),
         .M_Stage_sigma_constant_02_05(M_Stage_sigma_constant_02_05),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         M_Stage  me_14 (
         .out0(output_15_0),
         .in1(output_20_0),
         .in2(output_27_0),
         .in0(output_78_0),
         .in3(output_79_0),
         .M_Stage_sigma_constant_00_00(M_Stage_sigma_constant_00_00),
         .M_Stage_sigma_constant_01_01(M_Stage_sigma_constant_01_01),
         .M_Stage_sigma_constant_02_02(M_Stage_sigma_constant_02_02),
         .M_Stage_sigma_constant_00_03(M_Stage_sigma_constant_00_03),
         .M_Stage_sigma_constant_01_04(M_Stage_sigma_constant_01_04),
         .M_Stage_sigma_constant_02_05(M_Stage_sigma_constant_02_05),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         M_Stage  mf_15 (
         .out0(output_16_0),
         .in1(output_19_0),
         .in2(output_25_0),
         .in3(output_42_0),
         .in0(output_80_0),
         .M_Stage_sigma_constant_00_00(M_Stage_sigma_constant_00_00),
         .M_Stage_sigma_constant_01_01(M_Stage_sigma_constant_01_01),
         .M_Stage_sigma_constant_02_02(M_Stage_sigma_constant_02_02),
         .M_Stage_sigma_constant_00_03(M_Stage_sigma_constant_00_03),
         .M_Stage_sigma_constant_01_04(M_Stage_sigma_constant_01_04),
         .M_Stage_sigma_constant_02_05(M_Stage_sigma_constant_02_05),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Merge  merge_16 (
         .out0(output_17_0),
         .in0(output_1_0),
         .in1(output_2_0),
         .in2(output_3_0),
         .in3(output_4_0),
         .in4(output_5_0),
         .in5(output_6_0),
         .in6(output_7_0),
         .in7(output_8_0),
         .in8(output_9_0),
         .in9(output_10_0),
         .in10(output_11_0),
         .in11(output_12_0),
         .in12(output_13_0),
         .in13(output_14_0),
         .in14(output_15_0),
         .in15(output_16_0),
         .delay0(delay0),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer0_17 (
         .out0(output_19_0),
         .in0(output_14_0),
         .amount(M_buffer0_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer1_18 (
         .out0(output_20_0),
         .in0(output_13_0),
         .amount(M_buffer1_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer2_19 (
         .out0(output_21_0),
         .in0(output_12_0),
         .amount(M_buffer2_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer3_20 (
         .out0(output_22_0),
         .in0(output_11_0),
         .amount(M_buffer3_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer4_21 (
         .out0(output_23_0),
         .in0(output_10_0),
         .amount(M_buffer4_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer5_22 (
         .out0(output_24_0),
         .in0(output_9_0),
         .amount(M_buffer5_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer6_23 (
         .out0(output_25_0),
         .in0(output_9_0),
         .amount(M_buffer6_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer7_24 (
         .out0(output_26_0),
         .in0(output_8_0),
         .amount(M_buffer7_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer8_25 (
         .out0(output_27_0),
         .in0(output_8_0),
         .amount(M_buffer8_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer9_26 (
         .out0(output_28_0),
         .in0(output_7_0),
         .amount(M_buffer9_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer10_27 (
         .out0(output_29_0),
         .in0(output_7_0),
         .amount(M_buffer10_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer11_28 (
         .out0(output_30_0),
         .in0(output_6_0),
         .amount(M_buffer11_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer12_29 (
         .out0(output_31_0),
         .in0(output_6_0),
         .amount(M_buffer12_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer13_30 (
         .out0(output_32_0),
         .in0(output_5_0),
         .amount(M_buffer13_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer14_31 (
         .out0(output_33_0),
         .in0(output_5_0),
         .amount(M_buffer14_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer15_32 (
         .out0(output_34_0),
         .in0(output_4_0),
         .amount(M_buffer15_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer16_33 (
         .out0(output_35_0),
         .in0(output_4_0),
         .amount(M_buffer16_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer17_34 (
         .out0(output_36_0),
         .in0(output_3_0),
         .amount(M_buffer17_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer18_35 (
         .out0(output_37_0),
         .in0(output_3_0),
         .amount(M_buffer18_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer19_36 (
         .out0(output_38_0),
         .in0(output_2_0),
         .amount(M_buffer19_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer20_37 (
         .out0(output_39_0),
         .in0(output_2_0),
         .amount(M_buffer20_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer21_38 (
         .out0(output_40_0),
         .in0(output_1_0),
         .amount(M_buffer21_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer22_39 (
         .out0(output_41_0),
         .in0(output_1_0),
         .amount(M_buffer22_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer23_40 (
         .out0(output_42_0),
         .in0(output_1_0),
         .amount(M_buffer23_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer24_41 (
         .out0(output_43_0),
         .in0(in0), // w
         .amount(M_buffer24_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer25_42 (
         .out0(output_44_0),
         .in0(in0), // w
         .amount(M_buffer25_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer26_43 (
         .out0(output_45_0),
         .in0(in0), // w
         .amount(M_buffer26_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer27_44 (
         .out0(output_46_0),
         .in0(in0), // w
         .amount(M_buffer27_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer28_45 (
         .out0(output_47_0),
         .in0(in0), // w
         .amount(M_buffer28_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer29_46 (
         .out0(output_48_0),
         .in0(in0), // w
         .amount(M_buffer29_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer30_47 (
         .out0(output_49_0),
         .in0(in0), // w
         .amount(M_buffer30_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer31_48 (
         .out0(output_50_0),
         .in0(in0), // w
         .amount(M_buffer31_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer32_49 (
         .out0(output_51_0),
         .in0(in0), // w
         .amount(M_buffer32_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer33_50 (
         .out0(output_52_0),
         .in0(in0), // w
         .amount(M_buffer33_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer34_51 (
         .out0(output_53_0),
         .in0(in0), // w
         .amount(M_buffer34_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer35_52 (
         .out0(output_54_0),
         .in0(in0), // w
         .amount(M_buffer35_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer36_53 (
         .out0(output_55_0),
         .in0(in0), // w
         .amount(M_buffer36_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer37_54 (
         .out0(output_56_0),
         .in0(in0), // w
         .amount(M_buffer37_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer38_55 (
         .out0(output_57_0),
         .in0(in0), // w
         .amount(M_buffer38_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer39_56 (
         .out0(output_58_0),
         .in0(in0), // w
         .amount(M_buffer39_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer40_57 (
         .out0(output_59_0),
         .in0(in0), // w
         .amount(M_buffer40_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer41_58 (
         .out0(output_60_0),
         .in0(in0), // w
         .amount(M_buffer41_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer42_59 (
         .out0(output_61_0),
         .in0(in0), // w
         .amount(M_buffer42_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer43_60 (
         .out0(output_62_0),
         .in0(in0), // w
         .amount(M_buffer43_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer44_61 (
         .out0(output_63_0),
         .in0(in0), // w
         .amount(M_buffer44_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer45_62 (
         .out0(output_64_0),
         .in0(in0), // w
         .amount(M_buffer45_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer46_63 (
         .out0(output_65_0),
         .in0(in0), // w
         .amount(M_buffer46_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer47_64 (
         .out0(output_66_0),
         .in0(in0), // w
         .amount(M_buffer47_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer48_65 (
         .out0(output_67_0),
         .in0(in0), // w
         .amount(M_buffer48_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer49_66 (
         .out0(output_68_0),
         .in0(in0), // w
         .amount(M_buffer49_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer50_67 (
         .out0(output_69_0),
         .in0(in0), // w
         .amount(M_buffer50_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer51_68 (
         .out0(output_70_0),
         .in0(in0), // w
         .amount(M_buffer51_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer52_69 (
         .out0(output_71_0),
         .in0(in0), // w
         .amount(M_buffer52_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer53_70 (
         .out0(output_72_0),
         .in0(in0), // w
         .amount(M_buffer53_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer54_71 (
         .out0(output_73_0),
         .in0(in0), // w
         .amount(M_buffer54_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer55_72 (
         .out0(output_74_0),
         .in0(in0), // w
         .amount(M_buffer55_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer56_73 (
         .out0(output_75_0),
         .in0(in0), // w
         .amount(M_buffer56_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer57_74 (
         .out0(output_76_0),
         .in0(in0), // w
         .amount(M_buffer57_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer58_75 (
         .out0(output_77_0),
         .in0(in0), // w
         .amount(M_buffer58_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer59_76 (
         .out0(output_78_0),
         .in0(in0), // w
         .amount(M_buffer59_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer60_77 (
         .out0(output_79_0),
         .in0(in0), // w
         .amount(M_buffer60_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer61_78 (
         .out0(output_80_0),
         .in0(in0), // w
         .amount(M_buffer61_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         assign out0 = output_17_0;
   endmodule
