`timescale 1ns / 1ps
`include "global_defines.vh"
`include "system.vh"
`include "axi.vh"
`include "xversat.vh"
`include "xdefs.vh"

module ReadWriteAES #(
      parameter ADDR_W = `ADDR_W,
      parameter DATA_W = `DATA_W,
      parameter AXI_ADDR_W = 32
   )
   (

   input run,
   
   output done,
   input [31:0]     ext_addr_00,
   input [9:0]     int_addr_01,
   input [10:0]     size_02,
   input [9:0]     iterA_03,
   input [9:0]     perA_04,
   input [9:0]     dutyA_05,
   input [9:0]     shiftA_06,
   input [9:0]     incrA_07,
   input [7:0]     length_08,
   input [0:0]     pingPong_09,
   input [9:0]     iterB_10,
   input [9:0]     perB_11,
   input [9:0]     dutyB_12,
   input [9:0]     startB_13,
   input [9:0]     shiftB_14,
   input [9:0]     incrB_15,
   input [0:0]     reverseB_16,
   input [0:0]     extB_17,
   input [9:0]     iter2B_18,
   input [9:0]     per2B_19,
   input [9:0]     shift2B_20,
   input [9:0]     incr2B_21,
   input [31:0]     ext_addr_22,
   input [9:0]     int_addr_23,
   input [10:0]     size_24,
   input [9:0]     iterA_25,
   input [9:0]     perA_26,
   input [9:0]     dutyA_27,
   input [9:0]     shiftA_28,
   input [9:0]     incrA_29,
   input [7:0]     length_30,
   input [0:0]     pingPong_31,
   input [9:0]     iterB_32,
   input [9:0]     perB_33,
   input [9:0]     dutyB_34,
   input [9:0]     startB_35,
   input [9:0]     shiftB_36,
   input [9:0]     incrB_37,
   input [0:0]     reverseB_38,
   input [0:0]     extB_39,
   input [9:0]     iter2B_40,
   input [9:0]     per2B_41,
   input [9:0]     shift2B_42,
   input [9:0]     incr2B_43,
   input [31:0]     ext_addr_44,
   input [9:0]     int_addr_45,
   input [10:0]     size_46,
   input [9:0]     iterA_47,
   input [9:0]     perA_48,
   input [9:0]     dutyA_49,
   input [9:0]     shiftA_50,
   input [9:0]     incrA_51,
   input [7:0]     length_52,
   input [0:0]     pingPong_53,
   input [9:0]     iterB_54,
   input [9:0]     perB_55,
   input [9:0]     dutyB_56,
   input [9:0]     startB_57,
   input [9:0]     shiftB_58,
   input [9:0]     incrB_59,
   input [0:0]     reverseB_60,
   input [0:0]     extB_61,
   input [9:0]     iter2B_62,
   input [9:0]     per2B_63,
   input [9:0]     shift2B_64,
   input [9:0]     incr2B_65,
   input [31:0]     constant_00_66,
   input [31:0]     constant_01_67,
   input [31:0]     constant_02_68,
   input [31:0]     constant_03_69,
   input [31:0]     constant_04_70,
   input [31:0]     constant_05_71,
   input [31:0]     constant_06_72,
   input [31:0]     constant_07_73,
   input [31:0]     constant_08_74,
   input [31:0]     constant_09_75,
   input [5:0]     KeySchedule_buffer0_amount,
   input [5:0]     KeySchedule_buffer1_amount,
   input [5:0]     KeySchedule_buffer2_amount,
   input [5:0]     KeySchedule_buffer3_amount,
   input [5:0]     DoRow_buffer0_amount,
   input [5:0]     DoRow_buffer1_amount,
   input [5:0]     DoRow_buffer2_amount,
   input [5:0]     DoRow_buffer3_amount,
   input [5:0]     DoRow_buffer4_amount,
   input [5:0]     DoRow_buffer5_amount,
   input [5:0]     DoRow_buffer6_amount,
   input [5:0]     DoRow_buffer7_amount,
   input [5:0]     AES_buffer0_amount,
   input [5:0]     AES_buffer1_amount,
   input [5:0]     AES_buffer2_amount,
   input [5:0]     AES_buffer3_amount,
   input [5:0]     AES_buffer4_amount,
   input [5:0]     AES_buffer5_amount,
   input [5:0]     AES_buffer6_amount,
   input [5:0]     AES_buffer7_amount,
   input [5:0]     AES_buffer8_amount,
   input [5:0]     AES_buffer9_amount,
   input [5:0]     AES_buffer10_amount,
   input [5:0]     AES_buffer11_amount,
   input [5:0]     AES_buffer12_amount,
   input [5:0]     AES_buffer13_amount,
   input [5:0]     AES_buffer14_amount,
   input [5:0]     AES_buffer15_amount,
   input [5:0]     AES_buffer16_amount,
   input [5:0]     AES_buffer17_amount,
   input [5:0]     AES_buffer18_amount,
   input [5:0]     AES_buffer19_amount,
   input [5:0]     AES_buffer20_amount,
   input [5:0]     AES_buffer21_amount,
   input [5:0]     AES_buffer22_amount,
   input [5:0]     AES_buffer23_amount,
   input [5:0]     AES_buffer24_amount,
   input [5:0]     AES_buffer25_amount,
   input [5:0]     AES_buffer26_amount,
   input [5:0]     AES_buffer27_amount,
   input [5:0]     AES_buffer28_amount,
   input [5:0]     AES_buffer29_amount,
   input [5:0]     AES_buffer30_amount,
   input [5:0]     AES_buffer31_amount,
   input [5:0]     AES_buffer32_amount,
   input [5:0]     AES_buffer33_amount,
   input [5:0]     AES_buffer34_amount,
   input [5:0]     AES_buffer35_amount,
   input [5:0]     AES_buffer36_amount,
   input [5:0]     AES_buffer37_amount,
   input [5:0]     AES_buffer38_amount,
   input [5:0]     AES_buffer39_amount,
   input [5:0]     AES_buffer40_amount,
   input [5:0]     AES_buffer41_amount,
   input [5:0]     AES_buffer42_amount,
   input [5:0]     AES_buffer43_amount,
   input [5:0]     AES_buffer44_amount,
   input [5:0]     AES_buffer45_amount,
   input [5:0]     AES_buffer46_amount,
   input [5:0]     AES_buffer47_amount,
   input [5:0]     AES_buffer48_amount,
   input [5:0]     AES_buffer49_amount,
   input [5:0]     AES_buffer50_amount,
   input [5:0]     AES_buffer51_amount,
   input [5:0]     AES_buffer52_amount,
   input [5:0]     AES_buffer53_amount,
   input [5:0]     AES_buffer54_amount,
   input [5:0]     AES_buffer55_amount,
   input [5:0]     AES_buffer56_amount,
   input [5:0]     AES_buffer57_amount,
   input [5:0]     AES_buffer58_amount,
   input [5:0]     AES_buffer59_amount,
   input [5:0]     AES_buffer60_amount,
   input [5:0]     AES_buffer61_amount,
   input [5:0]     AES_buffer62_amount,
   input [5:0]     AES_buffer63_amount,
   input [5:0]     AES_buffer64_amount,
   input [5:0]     AES_buffer65_amount,
   input [5:0]     AES_buffer66_amount,
   input [5:0]     AES_buffer67_amount,
   input [5:0]     AES_buffer68_amount,
   input [5:0]     AES_buffer69_amount,
   input [5:0]     AES_buffer70_amount,
   input [5:0]     AES_buffer71_amount,
   input [5:0]     AES_buffer72_amount,
   input [5:0]     AES_buffer73_amount,
   input [5:0]     AES_buffer74_amount,
   input [5:0]     AES_buffer75_amount,
   input [5:0]     AES_buffer76_amount,
   input [5:0]     AES_buffer77_amount,
   input [5:0]     AES_buffer78_amount,
   input [5:0]     AES_buffer79_amount,
   input [5:0]     AES_buffer80_amount,
   input [5:0]     AES_buffer81_amount,
   input [5:0]     AES_buffer82_amount,
   input [5:0]     AES_buffer83_amount,
   input [5:0]     AES_buffer84_amount,
   input [5:0]     AES_buffer85_amount,
   input [5:0]     AES_buffer86_amount,
   input [5:0]     AES_buffer87_amount,
   input [5:0]     AES_buffer88_amount,
   input [5:0]     AES_buffer89_amount,
   input [5:0]     AES_buffer90_amount,
   input [5:0]     AES_buffer91_amount,
   input [5:0]     AES_buffer92_amount,
   input [5:0]     AES_buffer93_amount,
   input [5:0]     AES_buffer94_amount,
   input [5:0]     AES_buffer95_amount,
   input [5:0]     AES_buffer96_amount,
   input [5:0]     AES_buffer97_amount,
   input [5:0]     AES_buffer98_amount,
   input [5:0]     AES_buffer99_amount,
   input [5:0]     AES_buffer100_amount,
   input [5:0]     AES_buffer101_amount,
   input [5:0]     AES_buffer102_amount,
   input [5:0]     AES_buffer103_amount,
   input [5:0]     AES_buffer104_amount,
   input [5:0]     AES_buffer105_amount,
   input [5:0]     AES_buffer106_amount,
   input [5:0]     AES_buffer107_amount,
   input [5:0]     AES_buffer108_amount,
   input [5:0]     AES_buffer109_amount,
   input [5:0]     AES_buffer110_amount,
   input [5:0]     AES_buffer111_amount,
   input [5:0]     AES_buffer112_amount,
   input [5:0]     AES_buffer113_amount,
   input [5:0]     AES_buffer114_amount,
   input [5:0]     AES_buffer115_amount,
   input [5:0]     AES_buffer116_amount,
   input [5:0]     AES_buffer117_amount,
   input [5:0]     AES_buffer118_amount,
   input [5:0]     AES_buffer119_amount,
   input [5:0]     AES_buffer120_amount,
   input [5:0]     AES_buffer121_amount,
   input [5:0]     AES_buffer122_amount,
   input [5:0]     AES_buffer123_amount,
   input [5:0]     AES_buffer124_amount,
   input [5:0]     AES_buffer125_amount,
   input [5:0]     AES_buffer126_amount,
   input [5:0]     AES_buffer127_amount,
   input [5:0]     AES_buffer128_amount,
   input [5:0]     AES_buffer129_amount,
   input [5:0]     AES_buffer130_amount,
   input [5:0]     AES_buffer131_amount,
   input [5:0]     AES_buffer132_amount,
   input [5:0]     AES_buffer133_amount,
   input [5:0]     AES_buffer134_amount,
   input [5:0]     AES_buffer135_amount,
   input [5:0]     AES_buffer136_amount,
   input [5:0]     AES_buffer137_amount,
   input [5:0]     AES_buffer138_amount,
   input [5:0]     AES_buffer139_amount,
   input [5:0]     AES_buffer140_amount,
   input [5:0]     AES_buffer141_amount,
   input [5:0]     AES_buffer142_amount,
   input [5:0]     AES_buffer143_amount,
   input [5:0]     AES_buffer144_amount,
   input [5:0]     AES_buffer145_amount,
   input [5:0]     AES_buffer146_amount,
   input [5:0]     AES_buffer147_amount,
   input [5:0]     AES_buffer148_amount,
   input [5:0]     AES_buffer149_amount,
   input [5:0]     AES_buffer150_amount,
   input [5:0]     AES_buffer151_amount,
   input [5:0]     AES_buffer152_amount,
   input [5:0]     AES_buffer153_amount,
   input [5:0]     AES_buffer154_amount,
   input [5:0]     AES_buffer155_amount,
   input [5:0]     ReadWriteAES_buffer0_amount,
   input [5:0]     ReadWriteAES_buffer1_amount,
   input [5:0]     ReadWriteAES_buffer2_amount,
   input [5:0]     ReadWriteAES_buffer3_amount,
   input [5:0]     ReadWriteAES_buffer4_amount,
   input [5:0]     ReadWriteAES_buffer5_amount,
   input [5:0]     ReadWriteAES_buffer6_amount,
   input [5:0]     ReadWriteAES_buffer7_amount,
   input [5:0]     ReadWriteAES_buffer8_amount,
   input [5:0]     ReadWriteAES_buffer9_amount,
   input [5:0]     ReadWriteAES_buffer10_amount,
   input [5:0]     ReadWriteAES_buffer11_amount,
   input [5:0]     ReadWriteAES_buffer12_amount,
   input [5:0]     ReadWriteAES_buffer13_amount,
   input [5:0]     ReadWriteAES_buffer14_amount,
   input [5:0]     ReadWriteAES_buffer15_amount,
   input [5:0]     ReadWriteAES_buffer16_amount,
   input [5:0]     ReadWriteAES_buffer17_amount,
   input [5:0]     ReadWriteAES_buffer18_amount,
   input [5:0]     ReadWriteAES_buffer19_amount,
   input [5:0]     ReadWriteAES_buffer20_amount,
   input [5:0]     ReadWriteAES_buffer21_amount,
   input [5:0]     ReadWriteAES_buffer22_amount,
   input [5:0]     ReadWriteAES_buffer23_amount,
   input [5:0]     ReadWriteAES_buffer24_amount,
   input [5:0]     ReadWriteAES_buffer25_amount,
   input [5:0]     ReadWriteAES_buffer26_amount,
   input [5:0]     ReadWriteAES_buffer27_amount,
   input [5:0]     ReadWriteAES_buffer28_amount,
   input [5:0]     ReadWriteAES_buffer29_amount,
   input [5:0]     ReadWriteAES_buffer30_amount,
   input [5:0]     ReadWriteAES_buffer31_amount,
   input [5:0]     ReadWriteAES_buffer32_amount,
   input [5:0]     ReadWriteAES_buffer33_amount,
   input [5:0]     ReadWriteAES_buffer34_amount,
   input [5:0]     ReadWriteAES_buffer35_amount,
   input [5:0]     ReadWriteAES_buffer36_amount,
   input [5:0]     ReadWriteAES_buffer37_amount,
   input [5:0]     ReadWriteAES_buffer38_amount,
   input [5:0]     ReadWriteAES_buffer39_amount,
   input [5:0]     ReadWriteAES_buffer40_amount,
   input [5:0]     ReadWriteAES_buffer41_amount,
   input [5:0]     ReadWriteAES_buffer42_amount,
   input [5:0]     ReadWriteAES_buffer43_amount,
   input [5:0]     ReadWriteAES_buffer44_amount,
   input  [31:0]                   delay0,
   input  [31:0]                   delay1,
   input  [31:0]                   delay2,
   input  [31:0]                   delay3,
   // Databus master interface
   input [2:0]                databus_ready,
   output [2:0]               databus_valid,
   output [3 * AXI_ADDR_W-1:0]    databus_addr,
   input [`DATAPATH_W-1:0]                    databus_rdata,
   output [3 * `DATAPATH_W-1:0]   databus_wdata,
   output [3 * `DATAPATH_W/8-1:0] databus_wstrb,
   output [3 * 8-1:0]             databus_len,
   input  [2:0]               databus_last,
   // data/control interface
   input                           valid,
   input [16:0] addr,
   input [DATA_W/8-1:0]            wstrb,
   input [DATA_W-1:0]              wdata,
   output                          ready,
   output [DATA_W-1:0]             rdata,
   input                           clk,
   input                           rst
   );

wire wor_ready;

wire [31:0] unitRdataFinal;
reg [31:0] stateRead;

// Memory access
wire we = (|wstrb);
wire[0:0] unitReady;
reg [0:0] memoryMappedEnable;
wire [31:0] unitRData[0:0];

assign rdata = unitRdataFinal;
assign ready = wor_ready;
assign wor_ready = (|unitReady);

wire [31:0] rdata_0 ;

assign unitRdataFinal = (unitRData[0] );
wire [2:0] unitDone;
assign done = &unitDone;
wire [31:0] output_0_0 , output_1_0 , output_3_0 , output_4_0 , output_4_1 , output_4_2 , output_4_3 , output_4_4 , output_4_5 , output_4_6 , output_4_7 , output_4_8 , output_4_9 , output_4_10 , output_4_11 , output_4_12 , output_4_13 , output_4_14 , output_4_15 , output_5_0 , output_6_0 , output_7_0 , output_8_0 , output_9_0 , output_10_0 , output_11_0 , output_12_0 , output_13_0 , output_14_0 , output_15_0 , output_16_0 , output_17_0 , output_18_0 , output_19_0 , output_20_0 , output_21_0 , output_22_0 , output_23_0 , output_24_0 , output_25_0 , output_26_0 , output_27_0 , output_28_0 , output_29_0 , output_30_0 , output_31_0 , output_32_0 , output_33_0 , output_34_0 , output_35_0 , output_36_0 , output_37_0 , output_38_0 , output_39_0 , output_40_0 , output_41_0 , output_42_0 , output_43_0 , output_44_0 , output_45_0 , output_46_0 , output_47_0 , output_48_0 , output_49_0 ;

// Memory mapped
always @*
begin
   memoryMappedEnable = {1{1'b0}};
   if(valid)
   begin
   memoryMappedEnable[0] = 1'b1;
      end
end
VRead  cypher_0 (
         .out0(output_0_0),
         .ext_addr(ext_addr_00),
         .int_addr(int_addr_01),
         .size(size_02),
         .iterA(iterA_03),
         .perA(perA_04),
         .dutyA(dutyA_05),
         .shiftA(shiftA_06),
         .incrA(incrA_07),
         .length(length_08),
         .pingPong(pingPong_09),
         .iterB(iterB_10),
         .perB(perB_11),
         .dutyB(dutyB_12),
         .startB(startB_13),
         .shiftB(shiftB_14),
         .incrB(incrB_15),
         .reverseB(reverseB_16),
         .extB(extB_17),
         .iter2B(iter2B_18),
         .per2B(per2B_19),
         .shift2B(shift2B_20),
         .incr2B(incr2B_21),
         .delay0(delay0),
         .databus_ready(databus_ready[0 +: 1]),
         .databus_valid(databus_valid[0 +: 1]),
         .databus_addr(databus_addr[0 +: 32]),
         .databus_rdata(databus_rdata),
         .databus_wdata(databus_wdata[0 +: 32]),
         .databus_wstrb(databus_wstrb[0 +: 4]),
         .databus_len(databus_len[0 +: 8]),
         .databus_last(databus_last[0 +: 1]),
         .run(run),

         .done(unitDone[0]),
         .clk(clk),
         .rst(rst)
      );
         VRead  key_1 (
         .out0(output_1_0),
         .ext_addr(ext_addr_22),
         .int_addr(int_addr_23),
         .size(size_24),
         .iterA(iterA_25),
         .perA(perA_26),
         .dutyA(dutyA_27),
         .shiftA(shiftA_28),
         .incrA(incrA_29),
         .length(length_30),
         .pingPong(pingPong_31),
         .iterB(iterB_32),
         .perB(perB_33),
         .dutyB(dutyB_34),
         .startB(startB_35),
         .shiftB(shiftB_36),
         .incrB(incrB_37),
         .reverseB(reverseB_38),
         .extB(extB_39),
         .iter2B(iter2B_40),
         .per2B(per2B_41),
         .shift2B(shift2B_42),
         .incr2B(incr2B_43),
         .delay0(delay1),
         .databus_ready(databus_ready[1 +: 1]),
         .databus_valid(databus_valid[1 +: 1]),
         .databus_addr(databus_addr[32 +: 32]),
         .databus_rdata(databus_rdata),
         .databus_wdata(databus_wdata[32 +: 32]),
         .databus_wstrb(databus_wstrb[4 +: 4]),
         .databus_len(databus_len[8 +: 8]),
         .databus_last(databus_last[1 +: 1]),
         .run(run),

         .done(unitDone[1]),
         .clk(clk),
         .rst(rst)
      );
         VWrite  results_2 (
         .in0(output_3_0),
         .ext_addr(ext_addr_44),
         .int_addr(int_addr_45),
         .size(size_46),
         .iterA(iterA_47),
         .perA(perA_48),
         .dutyA(dutyA_49),
         .shiftA(shiftA_50),
         .incrA(incrA_51),
         .length(length_52),
         .pingPong(pingPong_53),
         .iterB(iterB_54),
         .perB(perB_55),
         .dutyB(dutyB_56),
         .startB(startB_57),
         .shiftB(shiftB_58),
         .incrB(incrB_59),
         .reverseB(reverseB_60),
         .extB(extB_61),
         .iter2B(iter2B_62),
         .per2B(per2B_63),
         .shift2B(shift2B_64),
         .incr2B(incr2B_65),
         .delay0(delay2),
         .databus_ready(databus_ready[2 +: 1]),
         .databus_valid(databus_valid[2 +: 1]),
         .databus_addr(databus_addr[64 +: 32]),
         .databus_rdata(databus_rdata),
         .databus_wdata(databus_wdata[64 +: 32]),
         .databus_wstrb(databus_wstrb[8 +: 4]),
         .databus_len(databus_len[16 +: 8]),
         .databus_last(databus_last[2 +: 1]),
         .run(run),

         .done(unitDone[2]),
         .clk(clk),
         .rst(rst)
      );
         Merge  merge_3 (
         .out0(output_3_0),
         .in0(output_4_0),
         .in1(output_5_0),
         .in2(output_6_0),
         .in3(output_7_0),
         .in4(output_8_0),
         .in5(output_9_0),
         .in6(output_10_0),
         .in7(output_11_0),
         .in8(output_12_0),
         .in9(output_13_0),
         .in10(output_14_0),
         .in11(output_15_0),
         .in12(output_16_0),
         .in13(output_17_0),
         .in14(output_18_0),
         .in15(output_19_0),
         .delay0(delay3),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         AES  aes_4 (
         .out0(output_4_0),
         .out1(output_4_1),
         .out2(output_4_2),
         .out3(output_4_3),
         .out4(output_4_4),
         .out5(output_4_5),
         .out6(output_4_6),
         .out7(output_4_7),
         .out8(output_4_8),
         .out9(output_4_9),
         .out10(output_4_10),
         .out11(output_4_11),
         .out12(output_4_12),
         .out13(output_4_13),
         .out14(output_4_14),
         .out15(output_4_15),
         .in15(output_0_0),
         .in31(output_1_0),
         .in16(output_20_0),
         .in17(output_21_0),
         .in18(output_22_0),
         .in19(output_23_0),
         .in20(output_24_0),
         .in21(output_25_0),
         .in22(output_26_0),
         .in23(output_27_0),
         .in24(output_28_0),
         .in25(output_29_0),
         .in26(output_30_0),
         .in27(output_31_0),
         .in28(output_32_0),
         .in29(output_33_0),
         .in30(output_34_0),
         .in0(output_35_0),
         .in1(output_36_0),
         .in2(output_37_0),
         .in3(output_38_0),
         .in4(output_39_0),
         .in5(output_40_0),
         .in6(output_41_0),
         .in7(output_42_0),
         .in8(output_43_0),
         .in9(output_44_0),
         .in10(output_45_0),
         .in11(output_46_0),
         .in12(output_47_0),
         .in13(output_48_0),
         .in14(output_49_0),
         .constant_00(constant_00_66),
         .constant_01(constant_01_67),
         .constant_02(constant_02_68),
         .constant_03(constant_03_69),
         .constant_04(constant_04_70),
         .constant_05(constant_05_71),
         .constant_06(constant_06_72),
         .constant_07(constant_07_73),
         .constant_08(constant_08_74),
         .constant_09(constant_09_75),
         .KeySchedule_buffer0_amount(KeySchedule_buffer0_amount),
         .KeySchedule_buffer1_amount(KeySchedule_buffer1_amount),
         .KeySchedule_buffer2_amount(KeySchedule_buffer2_amount),
         .KeySchedule_buffer3_amount(KeySchedule_buffer3_amount),
         .DoRow_buffer0_amount(DoRow_buffer0_amount),
         .DoRow_buffer1_amount(DoRow_buffer1_amount),
         .DoRow_buffer2_amount(DoRow_buffer2_amount),
         .DoRow_buffer3_amount(DoRow_buffer3_amount),
         .DoRow_buffer4_amount(DoRow_buffer4_amount),
         .DoRow_buffer5_amount(DoRow_buffer5_amount),
         .DoRow_buffer6_amount(DoRow_buffer6_amount),
         .DoRow_buffer7_amount(DoRow_buffer7_amount),
         .AES_buffer0_amount(AES_buffer0_amount),
         .AES_buffer1_amount(AES_buffer1_amount),
         .AES_buffer2_amount(AES_buffer2_amount),
         .AES_buffer3_amount(AES_buffer3_amount),
         .AES_buffer4_amount(AES_buffer4_amount),
         .AES_buffer5_amount(AES_buffer5_amount),
         .AES_buffer6_amount(AES_buffer6_amount),
         .AES_buffer7_amount(AES_buffer7_amount),
         .AES_buffer8_amount(AES_buffer8_amount),
         .AES_buffer9_amount(AES_buffer9_amount),
         .AES_buffer10_amount(AES_buffer10_amount),
         .AES_buffer11_amount(AES_buffer11_amount),
         .AES_buffer12_amount(AES_buffer12_amount),
         .AES_buffer13_amount(AES_buffer13_amount),
         .AES_buffer14_amount(AES_buffer14_amount),
         .AES_buffer15_amount(AES_buffer15_amount),
         .AES_buffer16_amount(AES_buffer16_amount),
         .AES_buffer17_amount(AES_buffer17_amount),
         .AES_buffer18_amount(AES_buffer18_amount),
         .AES_buffer19_amount(AES_buffer19_amount),
         .AES_buffer20_amount(AES_buffer20_amount),
         .AES_buffer21_amount(AES_buffer21_amount),
         .AES_buffer22_amount(AES_buffer22_amount),
         .AES_buffer23_amount(AES_buffer23_amount),
         .AES_buffer24_amount(AES_buffer24_amount),
         .AES_buffer25_amount(AES_buffer25_amount),
         .AES_buffer26_amount(AES_buffer26_amount),
         .AES_buffer27_amount(AES_buffer27_amount),
         .AES_buffer28_amount(AES_buffer28_amount),
         .AES_buffer29_amount(AES_buffer29_amount),
         .AES_buffer30_amount(AES_buffer30_amount),
         .AES_buffer31_amount(AES_buffer31_amount),
         .AES_buffer32_amount(AES_buffer32_amount),
         .AES_buffer33_amount(AES_buffer33_amount),
         .AES_buffer34_amount(AES_buffer34_amount),
         .AES_buffer35_amount(AES_buffer35_amount),
         .AES_buffer36_amount(AES_buffer36_amount),
         .AES_buffer37_amount(AES_buffer37_amount),
         .AES_buffer38_amount(AES_buffer38_amount),
         .AES_buffer39_amount(AES_buffer39_amount),
         .AES_buffer40_amount(AES_buffer40_amount),
         .AES_buffer41_amount(AES_buffer41_amount),
         .AES_buffer42_amount(AES_buffer42_amount),
         .AES_buffer43_amount(AES_buffer43_amount),
         .AES_buffer44_amount(AES_buffer44_amount),
         .AES_buffer45_amount(AES_buffer45_amount),
         .AES_buffer46_amount(AES_buffer46_amount),
         .AES_buffer47_amount(AES_buffer47_amount),
         .AES_buffer48_amount(AES_buffer48_amount),
         .AES_buffer49_amount(AES_buffer49_amount),
         .AES_buffer50_amount(AES_buffer50_amount),
         .AES_buffer51_amount(AES_buffer51_amount),
         .AES_buffer52_amount(AES_buffer52_amount),
         .AES_buffer53_amount(AES_buffer53_amount),
         .AES_buffer54_amount(AES_buffer54_amount),
         .AES_buffer55_amount(AES_buffer55_amount),
         .AES_buffer56_amount(AES_buffer56_amount),
         .AES_buffer57_amount(AES_buffer57_amount),
         .AES_buffer58_amount(AES_buffer58_amount),
         .AES_buffer59_amount(AES_buffer59_amount),
         .AES_buffer60_amount(AES_buffer60_amount),
         .AES_buffer61_amount(AES_buffer61_amount),
         .AES_buffer62_amount(AES_buffer62_amount),
         .AES_buffer63_amount(AES_buffer63_amount),
         .AES_buffer64_amount(AES_buffer64_amount),
         .AES_buffer65_amount(AES_buffer65_amount),
         .AES_buffer66_amount(AES_buffer66_amount),
         .AES_buffer67_amount(AES_buffer67_amount),
         .AES_buffer68_amount(AES_buffer68_amount),
         .AES_buffer69_amount(AES_buffer69_amount),
         .AES_buffer70_amount(AES_buffer70_amount),
         .AES_buffer71_amount(AES_buffer71_amount),
         .AES_buffer72_amount(AES_buffer72_amount),
         .AES_buffer73_amount(AES_buffer73_amount),
         .AES_buffer74_amount(AES_buffer74_amount),
         .AES_buffer75_amount(AES_buffer75_amount),
         .AES_buffer76_amount(AES_buffer76_amount),
         .AES_buffer77_amount(AES_buffer77_amount),
         .AES_buffer78_amount(AES_buffer78_amount),
         .AES_buffer79_amount(AES_buffer79_amount),
         .AES_buffer80_amount(AES_buffer80_amount),
         .AES_buffer81_amount(AES_buffer81_amount),
         .AES_buffer82_amount(AES_buffer82_amount),
         .AES_buffer83_amount(AES_buffer83_amount),
         .AES_buffer84_amount(AES_buffer84_amount),
         .AES_buffer85_amount(AES_buffer85_amount),
         .AES_buffer86_amount(AES_buffer86_amount),
         .AES_buffer87_amount(AES_buffer87_amount),
         .AES_buffer88_amount(AES_buffer88_amount),
         .AES_buffer89_amount(AES_buffer89_amount),
         .AES_buffer90_amount(AES_buffer90_amount),
         .AES_buffer91_amount(AES_buffer91_amount),
         .AES_buffer92_amount(AES_buffer92_amount),
         .AES_buffer93_amount(AES_buffer93_amount),
         .AES_buffer94_amount(AES_buffer94_amount),
         .AES_buffer95_amount(AES_buffer95_amount),
         .AES_buffer96_amount(AES_buffer96_amount),
         .AES_buffer97_amount(AES_buffer97_amount),
         .AES_buffer98_amount(AES_buffer98_amount),
         .AES_buffer99_amount(AES_buffer99_amount),
         .AES_buffer100_amount(AES_buffer100_amount),
         .AES_buffer101_amount(AES_buffer101_amount),
         .AES_buffer102_amount(AES_buffer102_amount),
         .AES_buffer103_amount(AES_buffer103_amount),
         .AES_buffer104_amount(AES_buffer104_amount),
         .AES_buffer105_amount(AES_buffer105_amount),
         .AES_buffer106_amount(AES_buffer106_amount),
         .AES_buffer107_amount(AES_buffer107_amount),
         .AES_buffer108_amount(AES_buffer108_amount),
         .AES_buffer109_amount(AES_buffer109_amount),
         .AES_buffer110_amount(AES_buffer110_amount),
         .AES_buffer111_amount(AES_buffer111_amount),
         .AES_buffer112_amount(AES_buffer112_amount),
         .AES_buffer113_amount(AES_buffer113_amount),
         .AES_buffer114_amount(AES_buffer114_amount),
         .AES_buffer115_amount(AES_buffer115_amount),
         .AES_buffer116_amount(AES_buffer116_amount),
         .AES_buffer117_amount(AES_buffer117_amount),
         .AES_buffer118_amount(AES_buffer118_amount),
         .AES_buffer119_amount(AES_buffer119_amount),
         .AES_buffer120_amount(AES_buffer120_amount),
         .AES_buffer121_amount(AES_buffer121_amount),
         .AES_buffer122_amount(AES_buffer122_amount),
         .AES_buffer123_amount(AES_buffer123_amount),
         .AES_buffer124_amount(AES_buffer124_amount),
         .AES_buffer125_amount(AES_buffer125_amount),
         .AES_buffer126_amount(AES_buffer126_amount),
         .AES_buffer127_amount(AES_buffer127_amount),
         .AES_buffer128_amount(AES_buffer128_amount),
         .AES_buffer129_amount(AES_buffer129_amount),
         .AES_buffer130_amount(AES_buffer130_amount),
         .AES_buffer131_amount(AES_buffer131_amount),
         .AES_buffer132_amount(AES_buffer132_amount),
         .AES_buffer133_amount(AES_buffer133_amount),
         .AES_buffer134_amount(AES_buffer134_amount),
         .AES_buffer135_amount(AES_buffer135_amount),
         .AES_buffer136_amount(AES_buffer136_amount),
         .AES_buffer137_amount(AES_buffer137_amount),
         .AES_buffer138_amount(AES_buffer138_amount),
         .AES_buffer139_amount(AES_buffer139_amount),
         .AES_buffer140_amount(AES_buffer140_amount),
         .AES_buffer141_amount(AES_buffer141_amount),
         .AES_buffer142_amount(AES_buffer142_amount),
         .AES_buffer143_amount(AES_buffer143_amount),
         .AES_buffer144_amount(AES_buffer144_amount),
         .AES_buffer145_amount(AES_buffer145_amount),
         .AES_buffer146_amount(AES_buffer146_amount),
         .AES_buffer147_amount(AES_buffer147_amount),
         .AES_buffer148_amount(AES_buffer148_amount),
         .AES_buffer149_amount(AES_buffer149_amount),
         .AES_buffer150_amount(AES_buffer150_amount),
         .AES_buffer151_amount(AES_buffer151_amount),
         .AES_buffer152_amount(AES_buffer152_amount),
         .AES_buffer153_amount(AES_buffer153_amount),
         .AES_buffer154_amount(AES_buffer154_amount),
         .AES_buffer155_amount(AES_buffer155_amount),
         .valid(memoryMappedEnable[0]),
         .wstrb(wstrb),
         .addr(addr[16:0]),
         .rdata(unitRData[0]),
         .ready(unitReady[0]),
         .wdata(wdata),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer0_5 (
         .out0(output_5_0),
         .in0(output_4_1),
         .amount(ReadWriteAES_buffer0_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer1_6 (
         .out0(output_6_0),
         .in0(output_4_2),
         .amount(ReadWriteAES_buffer1_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer2_7 (
         .out0(output_7_0),
         .in0(output_4_3),
         .amount(ReadWriteAES_buffer2_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer3_8 (
         .out0(output_8_0),
         .in0(output_4_4),
         .amount(ReadWriteAES_buffer3_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer4_9 (
         .out0(output_9_0),
         .in0(output_4_5),
         .amount(ReadWriteAES_buffer4_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer5_10 (
         .out0(output_10_0),
         .in0(output_4_6),
         .amount(ReadWriteAES_buffer5_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer6_11 (
         .out0(output_11_0),
         .in0(output_4_7),
         .amount(ReadWriteAES_buffer6_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer7_12 (
         .out0(output_12_0),
         .in0(output_4_8),
         .amount(ReadWriteAES_buffer7_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer8_13 (
         .out0(output_13_0),
         .in0(output_4_9),
         .amount(ReadWriteAES_buffer8_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer9_14 (
         .out0(output_14_0),
         .in0(output_4_10),
         .amount(ReadWriteAES_buffer9_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer10_15 (
         .out0(output_15_0),
         .in0(output_4_11),
         .amount(ReadWriteAES_buffer10_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer11_16 (
         .out0(output_16_0),
         .in0(output_4_12),
         .amount(ReadWriteAES_buffer11_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer12_17 (
         .out0(output_17_0),
         .in0(output_4_13),
         .amount(ReadWriteAES_buffer12_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer13_18 (
         .out0(output_18_0),
         .in0(output_4_14),
         .amount(ReadWriteAES_buffer13_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer14_19 (
         .out0(output_19_0),
         .in0(output_4_15),
         .amount(ReadWriteAES_buffer14_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer15_20 (
         .out0(output_20_0),
         .in0(output_1_0),
         .amount(ReadWriteAES_buffer15_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer16_21 (
         .out0(output_21_0),
         .in0(output_1_0),
         .amount(ReadWriteAES_buffer16_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer17_22 (
         .out0(output_22_0),
         .in0(output_1_0),
         .amount(ReadWriteAES_buffer17_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer18_23 (
         .out0(output_23_0),
         .in0(output_1_0),
         .amount(ReadWriteAES_buffer18_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer19_24 (
         .out0(output_24_0),
         .in0(output_1_0),
         .amount(ReadWriteAES_buffer19_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer20_25 (
         .out0(output_25_0),
         .in0(output_1_0),
         .amount(ReadWriteAES_buffer20_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer21_26 (
         .out0(output_26_0),
         .in0(output_1_0),
         .amount(ReadWriteAES_buffer21_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer22_27 (
         .out0(output_27_0),
         .in0(output_1_0),
         .amount(ReadWriteAES_buffer22_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer23_28 (
         .out0(output_28_0),
         .in0(output_1_0),
         .amount(ReadWriteAES_buffer23_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer24_29 (
         .out0(output_29_0),
         .in0(output_1_0),
         .amount(ReadWriteAES_buffer24_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer25_30 (
         .out0(output_30_0),
         .in0(output_1_0),
         .amount(ReadWriteAES_buffer25_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer26_31 (
         .out0(output_31_0),
         .in0(output_1_0),
         .amount(ReadWriteAES_buffer26_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer27_32 (
         .out0(output_32_0),
         .in0(output_1_0),
         .amount(ReadWriteAES_buffer27_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer28_33 (
         .out0(output_33_0),
         .in0(output_1_0),
         .amount(ReadWriteAES_buffer28_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer29_34 (
         .out0(output_34_0),
         .in0(output_1_0),
         .amount(ReadWriteAES_buffer29_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer30_35 (
         .out0(output_35_0),
         .in0(output_0_0),
         .amount(ReadWriteAES_buffer30_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer31_36 (
         .out0(output_36_0),
         .in0(output_0_0),
         .amount(ReadWriteAES_buffer31_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer32_37 (
         .out0(output_37_0),
         .in0(output_0_0),
         .amount(ReadWriteAES_buffer32_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer33_38 (
         .out0(output_38_0),
         .in0(output_0_0),
         .amount(ReadWriteAES_buffer33_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer34_39 (
         .out0(output_39_0),
         .in0(output_0_0),
         .amount(ReadWriteAES_buffer34_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer35_40 (
         .out0(output_40_0),
         .in0(output_0_0),
         .amount(ReadWriteAES_buffer35_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer36_41 (
         .out0(output_41_0),
         .in0(output_0_0),
         .amount(ReadWriteAES_buffer36_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer37_42 (
         .out0(output_42_0),
         .in0(output_0_0),
         .amount(ReadWriteAES_buffer37_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer38_43 (
         .out0(output_43_0),
         .in0(output_0_0),
         .amount(ReadWriteAES_buffer38_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer39_44 (
         .out0(output_44_0),
         .in0(output_0_0),
         .amount(ReadWriteAES_buffer39_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer40_45 (
         .out0(output_45_0),
         .in0(output_0_0),
         .amount(ReadWriteAES_buffer40_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer41_46 (
         .out0(output_46_0),
         .in0(output_0_0),
         .amount(ReadWriteAES_buffer41_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer42_47 (
         .out0(output_47_0),
         .in0(output_0_0),
         .amount(ReadWriteAES_buffer42_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer43_48 (
         .out0(output_48_0),
         .in0(output_0_0),
         .amount(ReadWriteAES_buffer43_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer44_49 (
         .out0(output_49_0),
         .in0(output_0_0),
         .amount(ReadWriteAES_buffer44_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         endmodule
