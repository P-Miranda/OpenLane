`define SRAM_ADDR_W 12
`define DATA_W 32
