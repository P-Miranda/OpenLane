`timescale 1ns / 1ps
`include "global_defines.vh"
`include "system.vh"
`include "axi.vh"
`include "xversat.vh"
`include "xdefs.vh"

module MatrixMultiplicationVread #(
      parameter ADDR_W = `ADDR_W,
      parameter DATA_W = `DATA_W,
      parameter AXI_ADDR_W = 32
   )
   (

   input run,
   
   output done,
   input [31:0]     ext_addr_00,
   input [9:0]     int_addr_01,
   input [10:0]     size_02,
   input [9:0]     iterA_03,
   input [9:0]     perA_04,
   input [9:0]     dutyA_05,
   input [9:0]     shiftA_06,
   input [9:0]     incrA_07,
   input [7:0]     length_08,
   input [0:0]     pingPong_09,
   input [9:0]     iterB_10,
   input [9:0]     perB_11,
   input [9:0]     dutyB_12,
   input [9:0]     startB_13,
   input [9:0]     shiftB_14,
   input [9:0]     incrB_15,
   input [0:0]     reverseB_16,
   input [0:0]     extB_17,
   input [9:0]     iter2B_18,
   input [9:0]     per2B_19,
   input [9:0]     shift2B_20,
   input [9:0]     incr2B_21,
   input [31:0]     ext_addr_22,
   input [9:0]     int_addr_23,
   input [10:0]     size_24,
   input [9:0]     iterA_25,
   input [9:0]     perA_26,
   input [9:0]     dutyA_27,
   input [9:0]     shiftA_28,
   input [9:0]     incrA_29,
   input [7:0]     length_30,
   input [0:0]     pingPong_31,
   input [9:0]     iterB_32,
   input [9:0]     perB_33,
   input [9:0]     dutyB_34,
   input [9:0]     startB_35,
   input [9:0]     shiftB_36,
   input [9:0]     incrB_37,
   input [0:0]     reverseB_38,
   input [0:0]     extB_39,
   input [9:0]     iter2B_40,
   input [9:0]     per2B_41,
   input [9:0]     shift2B_42,
   input [9:0]     incr2B_43,
   input [0:0]     opcode_44,
   input [9:0]     iterations_45,
   input [9:0]     period_46,
   input [5:0]     shift_47,
   input [31:0]     ext_addr_48,
   input [9:0]     int_addr_49,
   input [10:0]     size_50,
   input [9:0]     iterA_51,
   input [9:0]     perA_52,
   input [9:0]     dutyA_53,
   input [9:0]     shiftA_54,
   input [9:0]     incrA_55,
   input [7:0]     length_56,
   input [0:0]     pingPong_57,
   input [9:0]     iterB_58,
   input [9:0]     perB_59,
   input [9:0]     dutyB_60,
   input [9:0]     startB_61,
   input [9:0]     shiftB_62,
   input [9:0]     incrB_63,
   input [0:0]     reverseB_64,
   input [0:0]     extB_65,
   input [9:0]     iter2B_66,
   input [9:0]     per2B_67,
   input [9:0]     shift2B_68,
   input [9:0]     incr2B_69,
   input  [31:0]                   delay0,
   input  [31:0]                   delay1,
   input  [31:0]                   delay2,
   input  [31:0]                   delay3,
   // Databus master interface
   input [2:0]                databus_ready,
   output [2:0]               databus_valid,
   output [3 * AXI_ADDR_W-1:0]    databus_addr,
   input [`DATAPATH_W-1:0]                    databus_rdata,
   output [3 * `DATAPATH_W-1:0]   databus_wdata,
   output [3 * `DATAPATH_W/8-1:0] databus_wstrb,
   output [3 * 8-1:0]             databus_len,
   input  [2:0]               databus_last,
   input                           clk,
   input                           rst
   );

wire wor_ready;

wire [31:0] unitRdataFinal;
reg [31:0] stateRead;

wire [3:0] unitDone;
assign done = &unitDone;
wire [31:0] output_0_0 , output_1_0 , output_2_0 ;

VRead  matA_0 (
         .out0(output_0_0),
         .ext_addr(ext_addr_00),
         .int_addr(int_addr_01),
         .size(size_02),
         .iterA(iterA_03),
         .perA(perA_04),
         .dutyA(dutyA_05),
         .shiftA(shiftA_06),
         .incrA(incrA_07),
         .length(length_08),
         .pingPong(pingPong_09),
         .iterB(iterB_10),
         .perB(perB_11),
         .dutyB(dutyB_12),
         .startB(startB_13),
         .shiftB(shiftB_14),
         .incrB(incrB_15),
         .reverseB(reverseB_16),
         .extB(extB_17),
         .iter2B(iter2B_18),
         .per2B(per2B_19),
         .shift2B(shift2B_20),
         .incr2B(incr2B_21),
         .delay0(delay0),
         .databus_ready(databus_ready[0 +: 1]),
         .databus_valid(databus_valid[0 +: 1]),
         .databus_addr(databus_addr[0 +: 32]),
         .databus_rdata(databus_rdata),
         .databus_wdata(databus_wdata[0 +: 32]),
         .databus_wstrb(databus_wstrb[0 +: 4]),
         .databus_len(databus_len[0 +: 8]),
         .databus_last(databus_last[0 +: 1]),
         .run(run),

         .done(unitDone[0]),
         .clk(clk),
         .rst(rst)
      );
         VRead  matB_1 (
         .out0(output_1_0),
         .ext_addr(ext_addr_22),
         .int_addr(int_addr_23),
         .size(size_24),
         .iterA(iterA_25),
         .perA(perA_26),
         .dutyA(dutyA_27),
         .shiftA(shiftA_28),
         .incrA(incrA_29),
         .length(length_30),
         .pingPong(pingPong_31),
         .iterB(iterB_32),
         .perB(perB_33),
         .dutyB(dutyB_34),
         .startB(startB_35),
         .shiftB(shiftB_36),
         .incrB(incrB_37),
         .reverseB(reverseB_38),
         .extB(extB_39),
         .iter2B(iter2B_40),
         .per2B(per2B_41),
         .shift2B(shift2B_42),
         .incr2B(incr2B_43),
         .delay0(delay1),
         .databus_ready(databus_ready[1 +: 1]),
         .databus_valid(databus_valid[1 +: 1]),
         .databus_addr(databus_addr[32 +: 32]),
         .databus_rdata(databus_rdata),
         .databus_wdata(databus_wdata[32 +: 32]),
         .databus_wstrb(databus_wstrb[4 +: 4]),
         .databus_len(databus_len[8 +: 8]),
         .databus_last(databus_last[1 +: 1]),
         .run(run),

         .done(unitDone[1]),
         .clk(clk),
         .rst(rst)
      );
         Muladd  ma_2 (
         .out0(output_2_0),
         .in0(output_0_0),
         .in1(output_1_0),
         .opcode(opcode_44),
         .iterations(iterations_45),
         .period(period_46),
         .shift(shift_47),
         .delay0(delay2),
         .run(run),

         .done(unitDone[2]),
         .clk(clk),
         .rst(rst)
      );
         VWrite  res_3 (
         .in0(output_2_0),
         .ext_addr(ext_addr_48),
         .int_addr(int_addr_49),
         .size(size_50),
         .iterA(iterA_51),
         .perA(perA_52),
         .dutyA(dutyA_53),
         .shiftA(shiftA_54),
         .incrA(incrA_55),
         .length(length_56),
         .pingPong(pingPong_57),
         .iterB(iterB_58),
         .perB(perB_59),
         .dutyB(dutyB_60),
         .startB(startB_61),
         .shiftB(shiftB_62),
         .incrB(incrB_63),
         .reverseB(reverseB_64),
         .extB(extB_65),
         .iter2B(iter2B_66),
         .per2B(per2B_67),
         .shift2B(shift2B_68),
         .incr2B(incr2B_69),
         .delay0(delay3),
         .databus_ready(databus_ready[2 +: 1]),
         .databus_valid(databus_valid[2 +: 1]),
         .databus_addr(databus_addr[64 +: 32]),
         .databus_rdata(databus_rdata),
         .databus_wdata(databus_wdata[64 +: 32]),
         .databus_wstrb(databus_wstrb[8 +: 4]),
         .databus_len(databus_len[16 +: 8]),
         .databus_last(databus_last[2 +: 1]),
         .run(run),

         .done(unitDone[3]),
         .clk(clk),
         .rst(rst)
      );
         endmodule
