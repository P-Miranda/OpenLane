`define NUMBER_UNITS 1
`define CONFIG_W 1207
`define STATE_W 256
`define MAPPED_UNITS 1
`define MAPPED_BIT 13
`define nIO 1
`define VERSAT_IO
