`timescale 1ns / 1ps
`include "global_defines.vh"
`include "system.vh"
`include "axi.vh"
`include "xversat.vh"
`include "xdefs.vh"

module AES #(
      parameter ADDR_W = `ADDR_W,
      parameter DATA_W = `DATA_W,
      parameter AXI_ADDR_W = 32
   )
   (

   input run,
   
   input [DATA_W-1:0]              in0,
   input [DATA_W-1:0]              in1,
   input [DATA_W-1:0]              in2,
   input [DATA_W-1:0]              in3,
   input [DATA_W-1:0]              in4,
   input [DATA_W-1:0]              in5,
   input [DATA_W-1:0]              in6,
   input [DATA_W-1:0]              in7,
   input [DATA_W-1:0]              in8,
   input [DATA_W-1:0]              in9,
   input [DATA_W-1:0]              in10,
   input [DATA_W-1:0]              in11,
   input [DATA_W-1:0]              in12,
   input [DATA_W-1:0]              in13,
   input [DATA_W-1:0]              in14,
   input [DATA_W-1:0]              in15,
   input [DATA_W-1:0]              in16,
   input [DATA_W-1:0]              in17,
   input [DATA_W-1:0]              in18,
   input [DATA_W-1:0]              in19,
   input [DATA_W-1:0]              in20,
   input [DATA_W-1:0]              in21,
   input [DATA_W-1:0]              in22,
   input [DATA_W-1:0]              in23,
   input [DATA_W-1:0]              in24,
   input [DATA_W-1:0]              in25,
   input [DATA_W-1:0]              in26,
   input [DATA_W-1:0]              in27,
   input [DATA_W-1:0]              in28,
   input [DATA_W-1:0]              in29,
   input [DATA_W-1:0]              in30,
   input [DATA_W-1:0]              in31,
   output [DATA_W-1:0]             out0,
   output [DATA_W-1:0]             out1,
   output [DATA_W-1:0]             out2,
   output [DATA_W-1:0]             out3,
   output [DATA_W-1:0]             out4,
   output [DATA_W-1:0]             out5,
   output [DATA_W-1:0]             out6,
   output [DATA_W-1:0]             out7,
   output [DATA_W-1:0]             out8,
   output [DATA_W-1:0]             out9,
   output [DATA_W-1:0]             out10,
   output [DATA_W-1:0]             out11,
   output [DATA_W-1:0]             out12,
   output [DATA_W-1:0]             out13,
   output [DATA_W-1:0]             out14,
   output [DATA_W-1:0]             out15,
   input [31:0]     constant_00,
   input [31:0]     constant_01,
   input [31:0]     constant_02,
   input [31:0]     constant_03,
   input [31:0]     constant_04,
   input [31:0]     constant_05,
   input [31:0]     constant_06,
   input [31:0]     constant_07,
   input [31:0]     constant_08,
   input [31:0]     constant_09,
   input [5:0]     KeySchedule_buffer0_amount,
   input [5:0]     KeySchedule_buffer1_amount,
   input [5:0]     KeySchedule_buffer2_amount,
   input [5:0]     KeySchedule_buffer3_amount,
   input [5:0]     DoRow_buffer0_amount,
   input [5:0]     DoRow_buffer1_amount,
   input [5:0]     DoRow_buffer2_amount,
   input [5:0]     DoRow_buffer3_amount,
   input [5:0]     DoRow_buffer4_amount,
   input [5:0]     DoRow_buffer5_amount,
   input [5:0]     DoRow_buffer6_amount,
   input [5:0]     DoRow_buffer7_amount,
   input [5:0]     AES_buffer0_amount,
   input [5:0]     AES_buffer1_amount,
   input [5:0]     AES_buffer2_amount,
   input [5:0]     AES_buffer3_amount,
   input [5:0]     AES_buffer4_amount,
   input [5:0]     AES_buffer5_amount,
   input [5:0]     AES_buffer6_amount,
   input [5:0]     AES_buffer7_amount,
   input [5:0]     AES_buffer8_amount,
   input [5:0]     AES_buffer9_amount,
   input [5:0]     AES_buffer10_amount,
   input [5:0]     AES_buffer11_amount,
   input [5:0]     AES_buffer12_amount,
   input [5:0]     AES_buffer13_amount,
   input [5:0]     AES_buffer14_amount,
   input [5:0]     AES_buffer15_amount,
   input [5:0]     AES_buffer16_amount,
   input [5:0]     AES_buffer17_amount,
   input [5:0]     AES_buffer18_amount,
   input [5:0]     AES_buffer19_amount,
   input [5:0]     AES_buffer20_amount,
   input [5:0]     AES_buffer21_amount,
   input [5:0]     AES_buffer22_amount,
   input [5:0]     AES_buffer23_amount,
   input [5:0]     AES_buffer24_amount,
   input [5:0]     AES_buffer25_amount,
   input [5:0]     AES_buffer26_amount,
   input [5:0]     AES_buffer27_amount,
   input [5:0]     AES_buffer28_amount,
   input [5:0]     AES_buffer29_amount,
   input [5:0]     AES_buffer30_amount,
   input [5:0]     AES_buffer31_amount,
   input [5:0]     AES_buffer32_amount,
   input [5:0]     AES_buffer33_amount,
   input [5:0]     AES_buffer34_amount,
   input [5:0]     AES_buffer35_amount,
   input [5:0]     AES_buffer36_amount,
   input [5:0]     AES_buffer37_amount,
   input [5:0]     AES_buffer38_amount,
   input [5:0]     AES_buffer39_amount,
   input [5:0]     AES_buffer40_amount,
   input [5:0]     AES_buffer41_amount,
   input [5:0]     AES_buffer42_amount,
   input [5:0]     AES_buffer43_amount,
   input [5:0]     AES_buffer44_amount,
   input [5:0]     AES_buffer45_amount,
   input [5:0]     AES_buffer46_amount,
   input [5:0]     AES_buffer47_amount,
   input [5:0]     AES_buffer48_amount,
   input [5:0]     AES_buffer49_amount,
   input [5:0]     AES_buffer50_amount,
   input [5:0]     AES_buffer51_amount,
   input [5:0]     AES_buffer52_amount,
   input [5:0]     AES_buffer53_amount,
   input [5:0]     AES_buffer54_amount,
   input [5:0]     AES_buffer55_amount,
   input [5:0]     AES_buffer56_amount,
   input [5:0]     AES_buffer57_amount,
   input [5:0]     AES_buffer58_amount,
   input [5:0]     AES_buffer59_amount,
   input [5:0]     AES_buffer60_amount,
   input [5:0]     AES_buffer61_amount,
   input [5:0]     AES_buffer62_amount,
   input [5:0]     AES_buffer63_amount,
   input [5:0]     AES_buffer64_amount,
   input [5:0]     AES_buffer65_amount,
   input [5:0]     AES_buffer66_amount,
   input [5:0]     AES_buffer67_amount,
   input [5:0]     AES_buffer68_amount,
   input [5:0]     AES_buffer69_amount,
   input [5:0]     AES_buffer70_amount,
   input [5:0]     AES_buffer71_amount,
   input [5:0]     AES_buffer72_amount,
   input [5:0]     AES_buffer73_amount,
   input [5:0]     AES_buffer74_amount,
   input [5:0]     AES_buffer75_amount,
   input [5:0]     AES_buffer76_amount,
   input [5:0]     AES_buffer77_amount,
   input [5:0]     AES_buffer78_amount,
   input [5:0]     AES_buffer79_amount,
   input [5:0]     AES_buffer80_amount,
   input [5:0]     AES_buffer81_amount,
   input [5:0]     AES_buffer82_amount,
   input [5:0]     AES_buffer83_amount,
   input [5:0]     AES_buffer84_amount,
   input [5:0]     AES_buffer85_amount,
   input [5:0]     AES_buffer86_amount,
   input [5:0]     AES_buffer87_amount,
   input [5:0]     AES_buffer88_amount,
   input [5:0]     AES_buffer89_amount,
   input [5:0]     AES_buffer90_amount,
   input [5:0]     AES_buffer91_amount,
   input [5:0]     AES_buffer92_amount,
   input [5:0]     AES_buffer93_amount,
   input [5:0]     AES_buffer94_amount,
   input [5:0]     AES_buffer95_amount,
   input [5:0]     AES_buffer96_amount,
   input [5:0]     AES_buffer97_amount,
   input [5:0]     AES_buffer98_amount,
   input [5:0]     AES_buffer99_amount,
   input [5:0]     AES_buffer100_amount,
   input [5:0]     AES_buffer101_amount,
   input [5:0]     AES_buffer102_amount,
   input [5:0]     AES_buffer103_amount,
   input [5:0]     AES_buffer104_amount,
   input [5:0]     AES_buffer105_amount,
   input [5:0]     AES_buffer106_amount,
   input [5:0]     AES_buffer107_amount,
   input [5:0]     AES_buffer108_amount,
   input [5:0]     AES_buffer109_amount,
   input [5:0]     AES_buffer110_amount,
   input [5:0]     AES_buffer111_amount,
   input [5:0]     AES_buffer112_amount,
   input [5:0]     AES_buffer113_amount,
   input [5:0]     AES_buffer114_amount,
   input [5:0]     AES_buffer115_amount,
   input [5:0]     AES_buffer116_amount,
   input [5:0]     AES_buffer117_amount,
   input [5:0]     AES_buffer118_amount,
   input [5:0]     AES_buffer119_amount,
   input [5:0]     AES_buffer120_amount,
   input [5:0]     AES_buffer121_amount,
   input [5:0]     AES_buffer122_amount,
   input [5:0]     AES_buffer123_amount,
   input [5:0]     AES_buffer124_amount,
   input [5:0]     AES_buffer125_amount,
   input [5:0]     AES_buffer126_amount,
   input [5:0]     AES_buffer127_amount,
   input [5:0]     AES_buffer128_amount,
   input [5:0]     AES_buffer129_amount,
   input [5:0]     AES_buffer130_amount,
   input [5:0]     AES_buffer131_amount,
   input [5:0]     AES_buffer132_amount,
   input [5:0]     AES_buffer133_amount,
   input [5:0]     AES_buffer134_amount,
   input [5:0]     AES_buffer135_amount,
   input [5:0]     AES_buffer136_amount,
   input [5:0]     AES_buffer137_amount,
   input [5:0]     AES_buffer138_amount,
   input [5:0]     AES_buffer139_amount,
   input [5:0]     AES_buffer140_amount,
   input [5:0]     AES_buffer141_amount,
   input [5:0]     AES_buffer142_amount,
   input [5:0]     AES_buffer143_amount,
   input [5:0]     AES_buffer144_amount,
   input [5:0]     AES_buffer145_amount,
   input [5:0]     AES_buffer146_amount,
   input [5:0]     AES_buffer147_amount,
   input [5:0]     AES_buffer148_amount,
   input [5:0]     AES_buffer149_amount,
   input [5:0]     AES_buffer150_amount,
   input [5:0]     AES_buffer151_amount,
   input [5:0]     AES_buffer152_amount,
   input [5:0]     AES_buffer153_amount,
   input [5:0]     AES_buffer154_amount,
   input [5:0]     AES_buffer155_amount,
   // data/control interface
   input                           valid,
   input [16:0] addr,
   input [DATA_W/8-1:0]            wstrb,
   input [DATA_W-1:0]              wdata,
   output                          ready,
   output [DATA_W-1:0]             rdata,
   input                           clk,
   input                           rst
   );

wire wor_ready;

wire [31:0] unitRdataFinal;
reg [31:0] stateRead;

// Memory access
wire we = (|wstrb);
wire[19:0] unitReady;
reg [19:0] memoryMappedEnable;
wire [31:0] unitRData[19:0];

assign rdata = unitRdataFinal;
assign ready = wor_ready;
assign wor_ready = (|unitReady);

wire [31:0] rdata_0 , rdata_1 , rdata_2 , rdata_3 , rdata_4 , rdata_5 , rdata_6 , rdata_7 , rdata_8 , rdata_9 , rdata_10 , rdata_11 , rdata_12 , rdata_13 , rdata_14 , rdata_15 , rdata_16 , rdata_17 , rdata_18 , rdata_19 ;

assign unitRdataFinal = (unitRData[0] |unitRData[1] |unitRData[2] |unitRData[3] |unitRData[4] |unitRData[5] |unitRData[6] |unitRData[7] |unitRData[8] |unitRData[9] |unitRData[10] |unitRData[11] |unitRData[12] |unitRData[13] |unitRData[14] |unitRData[15] |unitRData[16] |unitRData[17] |unitRData[18] |unitRData[19] );
wire [31:0] output_0_0 , output_1_0 , output_2_0 , output_3_0 , output_4_0 , output_5_0 , output_6_0 , output_7_0 , output_8_0 , output_9_0 , output_10_0 , output_11_0 , output_12_0 , output_13_0 , output_14_0 , output_15_0 , output_16_0 , output_17_0 , output_18_0 , output_19_0 , output_20_0 , output_21_0 , output_22_0 , output_23_0 , output_24_0 , output_25_0 , output_26_0 , output_27_0 , output_28_0 , output_29_0 , output_30_0 , output_31_0 , output_32_0 , output_33_0 , output_34_0 , output_35_0 , output_36_0 , output_37_0 , output_38_0 , output_39_0 , output_40_0 , output_41_0 , output_42_0 , output_42_1 , output_42_2 , output_42_3 , output_42_4 , output_42_5 , output_42_6 , output_42_7 , output_42_8 , output_42_9 , output_42_10 , output_42_11 , output_42_12 , output_42_13 , output_42_14 , output_42_15 , output_43_0 , output_43_1 , output_43_2 , output_43_3 , output_43_4 , output_43_5 , output_43_6 , output_43_7 , output_43_8 , output_43_9 , output_43_10 , output_43_11 , output_43_12 , output_43_13 , output_43_14 , output_43_15 , output_44_0 , output_44_1 , output_44_2 , output_44_3 , output_44_4 , output_44_5 , output_44_6 , output_44_7 , output_44_8 , output_44_9 , output_44_10 , output_44_11 , output_44_12 , output_44_13 , output_44_14 , output_44_15 , output_45_0 , output_45_1 , output_45_2 , output_45_3 , output_45_4 , output_45_5 , output_45_6 , output_45_7 , output_45_8 , output_45_9 , output_45_10 , output_45_11 , output_45_12 , output_45_13 , output_45_14 , output_45_15 , output_46_0 , output_46_1 , output_46_2 , output_46_3 , output_46_4 , output_46_5 , output_46_6 , output_46_7 , output_46_8 , output_46_9 , output_46_10 , output_46_11 , output_46_12 , output_46_13 , output_46_14 , output_46_15 , output_47_0 , output_47_1 , output_47_2 , output_47_3 , output_47_4 , output_47_5 , output_47_6 , output_47_7 , output_47_8 , output_47_9 , output_47_10 , output_47_11 , output_47_12 , output_47_13 , output_47_14 , output_47_15 , output_48_0 , output_48_1 , output_48_2 , output_48_3 , output_48_4 , output_48_5 , output_48_6 , output_48_7 , output_48_8 , output_48_9 , output_48_10 , output_48_11 , output_48_12 , output_48_13 , output_48_14 , output_48_15 , output_49_0 , output_49_1 , output_49_2 , output_49_3 , output_49_4 , output_49_5 , output_49_6 , output_49_7 , output_49_8 , output_49_9 , output_49_10 , output_49_11 , output_49_12 , output_49_13 , output_49_14 , output_49_15 , output_50_0 , output_50_1 , output_50_2 , output_50_3 , output_50_4 , output_50_5 , output_50_6 , output_50_7 , output_50_8 , output_50_9 , output_50_10 , output_50_11 , output_50_12 , output_50_13 , output_50_14 , output_50_15 , output_51_0 , output_51_1 , output_51_2 , output_51_3 , output_51_4 , output_51_5 , output_51_6 , output_51_7 , output_51_8 , output_51_9 , output_51_10 , output_51_11 , output_51_12 , output_51_13 , output_51_14 , output_51_15 , output_52_0 , output_52_1 , output_52_2 , output_52_3 , output_52_4 , output_52_5 , output_52_6 , output_52_7 , output_52_8 , output_52_9 , output_52_10 , output_52_11 , output_52_12 , output_52_13 , output_52_14 , output_52_15 , output_53_0 , output_53_1 , output_53_2 , output_53_3 , output_53_4 , output_53_5 , output_53_6 , output_53_7 , output_53_8 , output_53_9 , output_53_10 , output_53_11 , output_53_12 , output_53_13 , output_53_14 , output_53_15 , output_54_0 , output_54_1 , output_54_2 , output_54_3 , output_54_4 , output_54_5 , output_54_6 , output_54_7 , output_54_8 , output_54_9 , output_54_10 , output_54_11 , output_54_12 , output_54_13 , output_54_14 , output_54_15 , output_55_0 , output_55_1 , output_55_2 , output_55_3 , output_55_4 , output_55_5 , output_55_6 , output_55_7 , output_55_8 , output_55_9 , output_55_10 , output_55_11 , output_55_12 , output_55_13 , output_55_14 , output_55_15 , output_56_0 , output_56_1 , output_56_2 , output_56_3 , output_56_4 , output_56_5 , output_56_6 , output_56_7 , output_56_8 , output_56_9 , output_56_10 , output_56_11 , output_56_12 , output_56_13 , output_56_14 , output_56_15 , output_57_0 , output_57_1 , output_57_2 , output_57_3 , output_57_4 , output_57_5 , output_57_6 , output_57_7 , output_57_8 , output_57_9 , output_57_10 , output_57_11 , output_57_12 , output_57_13 , output_57_14 , output_57_15 , output_58_0 , output_58_1 , output_58_2 , output_58_3 , output_58_4 , output_58_5 , output_58_6 , output_58_7 , output_58_8 , output_58_9 , output_58_10 , output_58_11 , output_58_12 , output_58_13 , output_58_14 , output_58_15 , output_59_0 , output_59_1 , output_59_2 , output_59_3 , output_59_4 , output_59_5 , output_59_6 , output_59_7 , output_59_8 , output_59_9 , output_59_10 , output_59_11 , output_59_12 , output_59_13 , output_59_14 , output_59_15 , output_60_0 , output_60_1 , output_60_2 , output_60_3 , output_60_4 , output_60_5 , output_60_6 , output_60_7 , output_60_8 , output_60_9 , output_60_10 , output_60_11 , output_60_12 , output_60_13 , output_60_14 , output_60_15 , output_61_0 , output_61_1 , output_61_2 , output_61_3 , output_61_4 , output_61_5 , output_61_6 , output_61_7 , output_61_8 , output_61_9 , output_61_10 , output_61_11 , output_61_12 , output_61_13 , output_61_14 , output_61_15 , output_62_0 , output_62_1 , output_62_2 , output_62_3 , output_62_4 , output_62_5 , output_62_6 , output_62_7 , output_62_8 , output_62_9 , output_62_10 , output_62_11 , output_62_12 , output_62_13 , output_62_14 , output_62_15 , output_63_0 , output_63_1 , output_63_2 , output_63_3 , output_63_4 , output_63_5 , output_63_6 , output_63_7 , output_63_8 , output_63_9 , output_63_10 , output_63_11 , output_63_12 , output_63_13 , output_63_14 , output_63_15 , output_64_0 , output_64_1 , output_64_2 , output_64_3 , output_64_4 , output_64_5 , output_64_6 , output_64_7 , output_64_8 , output_64_9 , output_64_10 , output_64_11 , output_64_12 , output_64_13 , output_64_14 , output_64_15 , output_66_0 , output_67_0 , output_68_0 , output_69_0 , output_70_0 , output_71_0 , output_72_0 , output_73_0 , output_74_0 , output_75_0 , output_76_0 , output_77_0 , output_78_0 , output_79_0 , output_80_0 , output_81_0 , output_82_0 , output_83_0 , output_84_0 , output_85_0 , output_86_0 , output_87_0 , output_88_0 , output_89_0 , output_90_0 , output_91_0 , output_92_0 , output_93_0 , output_94_0 , output_95_0 , output_96_0 , output_97_0 , output_98_0 , output_99_0 , output_100_0 , output_101_0 , output_102_0 , output_103_0 , output_104_0 , output_105_0 , output_106_0 , output_107_0 , output_108_0 , output_109_0 , output_110_0 , output_111_0 , output_112_0 , output_113_0 , output_114_0 , output_115_0 , output_116_0 , output_117_0 , output_118_0 , output_119_0 , output_120_0 , output_121_0 , output_122_0 , output_123_0 , output_124_0 , output_125_0 , output_126_0 , output_127_0 , output_128_0 , output_129_0 , output_130_0 , output_131_0 , output_132_0 , output_133_0 , output_134_0 , output_135_0 , output_136_0 , output_137_0 , output_138_0 , output_139_0 , output_140_0 , output_141_0 , output_142_0 , output_143_0 , output_144_0 , output_145_0 , output_146_0 , output_147_0 , output_148_0 , output_149_0 , output_150_0 , output_151_0 , output_152_0 , output_153_0 , output_154_0 , output_155_0 , output_156_0 , output_157_0 , output_158_0 , output_159_0 , output_160_0 , output_161_0 , output_162_0 , output_163_0 , output_164_0 , output_165_0 , output_166_0 , output_167_0 , output_168_0 , output_169_0 , output_170_0 , output_171_0 , output_172_0 , output_173_0 , output_174_0 , output_175_0 , output_176_0 , output_177_0 , output_178_0 , output_179_0 , output_180_0 , output_181_0 , output_182_0 , output_183_0 , output_184_0 , output_185_0 , output_186_0 , output_187_0 , output_188_0 , output_189_0 , output_190_0 , output_191_0 , output_192_0 , output_193_0 , output_194_0 , output_195_0 , output_196_0 , output_197_0 , output_198_0 , output_199_0 , output_200_0 , output_201_0 , output_202_0 , output_203_0 , output_204_0 , output_205_0 , output_206_0 , output_207_0 , output_208_0 , output_209_0 , output_210_0 , output_211_0 , output_212_0 , output_213_0 , output_214_0 , output_215_0 , output_216_0 , output_217_0 , output_218_0 , output_219_0 , output_220_0 , output_221_0 ;

// Memory mapped
always @*
begin
   memoryMappedEnable = {20{1'b0}};
   if(valid)
   begin
   if(addr[16:9] == 8'b00100111)
            memoryMappedEnable[0] = 1'b1;
      if(addr[16:9] == 8'b00100001)
            memoryMappedEnable[1] = 1'b1;
      if(addr[16:9] == 8'b00100110)
            memoryMappedEnable[2] = 1'b1;
      if(addr[16:10] == 7'b0010110)
            memoryMappedEnable[3] = 1'b1;
      if(addr[16:9] == 8'b00100000)
            memoryMappedEnable[4] = 1'b1;
      if(addr[16:9] == 8'b00100010)
            memoryMappedEnable[5] = 1'b1;
      if(addr[16:9] == 8'b00100011)
            memoryMappedEnable[6] = 1'b1;
      if(addr[16:9] == 8'b00100100)
            memoryMappedEnable[7] = 1'b1;
      if(addr[16:9] == 8'b00100101)
            memoryMappedEnable[8] = 1'b1;
      if(addr[16:10] == 7'b0010111)
            memoryMappedEnable[9] = 1'b1;
      if(addr[16:13] == 4'b0000)
            memoryMappedEnable[10] = 1'b1;
      if(addr[16:14] == 3'b010)
            memoryMappedEnable[11] = 1'b1;
      if(addr[16:14] == 3'b101)
            memoryMappedEnable[12] = 1'b1;
      if(addr[16:13] == 4'b0001)
            memoryMappedEnable[13] = 1'b1;
      if(addr[16:14] == 3'b011)
            memoryMappedEnable[14] = 1'b1;
      if(addr[16:13] == 4'b0011)
            memoryMappedEnable[15] = 1'b1;
      if(addr[16:14] == 3'b110)
            memoryMappedEnable[16] = 1'b1;
      if(addr[16:14] == 3'b111)
            memoryMappedEnable[17] = 1'b1;
      if(addr[16:14] == 3'b100)
            memoryMappedEnable[18] = 1'b1;
      if(addr[16:11] == 6'b001010)
            memoryMappedEnable[19] = 1'b1;
      end
end
Const  rcon0_0 (
         .out0(output_32_0),
         .constant(constant_00),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Const  rcon1_1 (
         .out0(output_33_0),
         .constant(constant_01),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Const  rcon2_2 (
         .out0(output_34_0),
         .constant(constant_02),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Const  rcon3_3 (
         .out0(output_35_0),
         .constant(constant_03),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Const  rcon4_4 (
         .out0(output_36_0),
         .constant(constant_04),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Const  rcon5_5 (
         .out0(output_37_0),
         .constant(constant_05),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Const  rcon6_6 (
         .out0(output_38_0),
         .constant(constant_06),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Const  rcon7_7 (
         .out0(output_39_0),
         .constant(constant_07),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Const  rcon8_8 (
         .out0(output_40_0),
         .constant(constant_08),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Const  rcon9_9 (
         .out0(output_41_0),
         .constant(constant_09),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         KeySchedule  key0_10 (
         .out0(output_42_0),
         .out1(output_42_1),
         .out2(output_42_2),
         .out3(output_42_3),
         .out4(output_42_4),
         .out5(output_42_5),
         .out6(output_42_6),
         .out7(output_42_7),
         .out8(output_42_8),
         .out9(output_42_9),
         .out10(output_42_10),
         .out11(output_42_11),
         .out12(output_42_12),
         .out13(output_42_13),
         .out14(output_42_14),
         .out15(output_42_15),
         .in16(output_32_0),
         .in15(output_206_0),
         .in14(output_207_0),
         .in13(output_208_0),
         .in12(output_209_0),
         .in11(output_210_0),
         .in10(output_211_0),
         .in9(output_212_0),
         .in8(output_213_0),
         .in7(output_214_0),
         .in6(output_215_0),
         .in5(output_216_0),
         .in4(output_217_0),
         .in3(output_218_0),
         .in2(output_219_0),
         .in1(output_220_0),
         .in0(output_221_0),
         .KeySchedule_buffer0_amount(KeySchedule_buffer0_amount),
         .KeySchedule_buffer1_amount(KeySchedule_buffer1_amount),
         .KeySchedule_buffer2_amount(KeySchedule_buffer2_amount),
         .KeySchedule_buffer3_amount(KeySchedule_buffer3_amount),
         .valid(memoryMappedEnable[0]),
         .wstrb(wstrb),
         .addr(addr[8:0]),
         .rdata(unitRData[0]),
         .ready(unitReady[0]),
         .wdata(wdata),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         KeySchedule  key1_11 (
         .out0(output_43_0),
         .out1(output_43_1),
         .out2(output_43_2),
         .out3(output_43_3),
         .out4(output_43_4),
         .out5(output_43_5),
         .out6(output_43_6),
         .out7(output_43_7),
         .out8(output_43_8),
         .out9(output_43_9),
         .out10(output_43_10),
         .out11(output_43_11),
         .out12(output_43_12),
         .out13(output_43_13),
         .out14(output_43_14),
         .out15(output_43_15),
         .in16(output_33_0),
         .in0(output_190_0),
         .in1(output_191_0),
         .in2(output_192_0),
         .in3(output_193_0),
         .in4(output_194_0),
         .in5(output_195_0),
         .in6(output_196_0),
         .in7(output_197_0),
         .in8(output_198_0),
         .in9(output_199_0),
         .in10(output_200_0),
         .in11(output_201_0),
         .in12(output_202_0),
         .in13(output_203_0),
         .in14(output_204_0),
         .in15(output_205_0),
         .KeySchedule_buffer0_amount(KeySchedule_buffer0_amount),
         .KeySchedule_buffer1_amount(KeySchedule_buffer1_amount),
         .KeySchedule_buffer2_amount(KeySchedule_buffer2_amount),
         .KeySchedule_buffer3_amount(KeySchedule_buffer3_amount),
         .valid(memoryMappedEnable[1]),
         .wstrb(wstrb),
         .addr(addr[8:0]),
         .rdata(unitRData[1]),
         .ready(unitReady[1]),
         .wdata(wdata),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         KeySchedule  key2_12 (
         .out0(output_44_0),
         .out1(output_44_1),
         .out2(output_44_2),
         .out3(output_44_3),
         .out4(output_44_4),
         .out5(output_44_5),
         .out6(output_44_6),
         .out7(output_44_7),
         .out8(output_44_8),
         .out9(output_44_9),
         .out10(output_44_10),
         .out11(output_44_11),
         .out12(output_44_12),
         .out13(output_44_13),
         .out14(output_44_14),
         .out15(output_44_15),
         .in16(output_34_0),
         .in0(output_174_0),
         .in1(output_175_0),
         .in2(output_176_0),
         .in3(output_177_0),
         .in4(output_178_0),
         .in5(output_179_0),
         .in6(output_180_0),
         .in7(output_181_0),
         .in8(output_182_0),
         .in9(output_183_0),
         .in10(output_184_0),
         .in11(output_185_0),
         .in12(output_186_0),
         .in13(output_187_0),
         .in14(output_188_0),
         .in15(output_189_0),
         .KeySchedule_buffer0_amount(KeySchedule_buffer0_amount),
         .KeySchedule_buffer1_amount(KeySchedule_buffer1_amount),
         .KeySchedule_buffer2_amount(KeySchedule_buffer2_amount),
         .KeySchedule_buffer3_amount(KeySchedule_buffer3_amount),
         .valid(memoryMappedEnable[2]),
         .wstrb(wstrb),
         .addr(addr[8:0]),
         .rdata(unitRData[2]),
         .ready(unitReady[2]),
         .wdata(wdata),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         KeySchedule  key3_13 (
         .out0(output_45_0),
         .out1(output_45_1),
         .out2(output_45_2),
         .out3(output_45_3),
         .out4(output_45_4),
         .out5(output_45_5),
         .out6(output_45_6),
         .out7(output_45_7),
         .out8(output_45_8),
         .out9(output_45_9),
         .out10(output_45_10),
         .out11(output_45_11),
         .out12(output_45_12),
         .out13(output_45_13),
         .out14(output_45_14),
         .out15(output_45_15),
         .in16(output_35_0),
         .in0(output_158_0),
         .in1(output_159_0),
         .in2(output_160_0),
         .in3(output_161_0),
         .in4(output_162_0),
         .in5(output_163_0),
         .in6(output_164_0),
         .in7(output_165_0),
         .in8(output_166_0),
         .in9(output_167_0),
         .in10(output_168_0),
         .in11(output_169_0),
         .in12(output_170_0),
         .in13(output_171_0),
         .in14(output_172_0),
         .in15(output_173_0),
         .KeySchedule_buffer0_amount(KeySchedule_buffer0_amount),
         .KeySchedule_buffer1_amount(KeySchedule_buffer1_amount),
         .KeySchedule_buffer2_amount(KeySchedule_buffer2_amount),
         .KeySchedule_buffer3_amount(KeySchedule_buffer3_amount),
         .valid(memoryMappedEnable[3]),
         .wstrb(wstrb),
         .addr(addr[8:0]),
         .rdata(unitRData[3]),
         .ready(unitReady[3]),
         .wdata(wdata),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         KeySchedule  key4_14 (
         .out0(output_46_0),
         .out1(output_46_1),
         .out2(output_46_2),
         .out3(output_46_3),
         .out4(output_46_4),
         .out5(output_46_5),
         .out6(output_46_6),
         .out7(output_46_7),
         .out8(output_46_8),
         .out9(output_46_9),
         .out10(output_46_10),
         .out11(output_46_11),
         .out12(output_46_12),
         .out13(output_46_13),
         .out14(output_46_14),
         .out15(output_46_15),
         .in16(output_36_0),
         .in0(output_142_0),
         .in1(output_143_0),
         .in2(output_144_0),
         .in3(output_145_0),
         .in4(output_146_0),
         .in5(output_147_0),
         .in6(output_148_0),
         .in7(output_149_0),
         .in8(output_150_0),
         .in9(output_151_0),
         .in10(output_152_0),
         .in11(output_153_0),
         .in12(output_154_0),
         .in13(output_155_0),
         .in14(output_156_0),
         .in15(output_157_0),
         .KeySchedule_buffer0_amount(KeySchedule_buffer0_amount),
         .KeySchedule_buffer1_amount(KeySchedule_buffer1_amount),
         .KeySchedule_buffer2_amount(KeySchedule_buffer2_amount),
         .KeySchedule_buffer3_amount(KeySchedule_buffer3_amount),
         .valid(memoryMappedEnable[4]),
         .wstrb(wstrb),
         .addr(addr[8:0]),
         .rdata(unitRData[4]),
         .ready(unitReady[4]),
         .wdata(wdata),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         KeySchedule  key5_15 (
         .out0(output_47_0),
         .out1(output_47_1),
         .out2(output_47_2),
         .out3(output_47_3),
         .out4(output_47_4),
         .out5(output_47_5),
         .out6(output_47_6),
         .out7(output_47_7),
         .out8(output_47_8),
         .out9(output_47_9),
         .out10(output_47_10),
         .out11(output_47_11),
         .out12(output_47_12),
         .out13(output_47_13),
         .out14(output_47_14),
         .out15(output_47_15),
         .in16(output_37_0),
         .in0(output_126_0),
         .in1(output_127_0),
         .in2(output_128_0),
         .in3(output_129_0),
         .in4(output_130_0),
         .in5(output_131_0),
         .in6(output_132_0),
         .in7(output_133_0),
         .in8(output_134_0),
         .in9(output_135_0),
         .in10(output_136_0),
         .in11(output_137_0),
         .in12(output_138_0),
         .in13(output_139_0),
         .in14(output_140_0),
         .in15(output_141_0),
         .KeySchedule_buffer0_amount(KeySchedule_buffer0_amount),
         .KeySchedule_buffer1_amount(KeySchedule_buffer1_amount),
         .KeySchedule_buffer2_amount(KeySchedule_buffer2_amount),
         .KeySchedule_buffer3_amount(KeySchedule_buffer3_amount),
         .valid(memoryMappedEnable[5]),
         .wstrb(wstrb),
         .addr(addr[8:0]),
         .rdata(unitRData[5]),
         .ready(unitReady[5]),
         .wdata(wdata),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         KeySchedule  key6_16 (
         .out0(output_48_0),
         .out1(output_48_1),
         .out2(output_48_2),
         .out3(output_48_3),
         .out4(output_48_4),
         .out5(output_48_5),
         .out6(output_48_6),
         .out7(output_48_7),
         .out8(output_48_8),
         .out9(output_48_9),
         .out10(output_48_10),
         .out11(output_48_11),
         .out12(output_48_12),
         .out13(output_48_13),
         .out14(output_48_14),
         .out15(output_48_15),
         .in16(output_38_0),
         .in0(output_110_0),
         .in1(output_111_0),
         .in2(output_112_0),
         .in3(output_113_0),
         .in4(output_114_0),
         .in5(output_115_0),
         .in6(output_116_0),
         .in7(output_117_0),
         .in8(output_118_0),
         .in9(output_119_0),
         .in10(output_120_0),
         .in11(output_121_0),
         .in12(output_122_0),
         .in13(output_123_0),
         .in14(output_124_0),
         .in15(output_125_0),
         .KeySchedule_buffer0_amount(KeySchedule_buffer0_amount),
         .KeySchedule_buffer1_amount(KeySchedule_buffer1_amount),
         .KeySchedule_buffer2_amount(KeySchedule_buffer2_amount),
         .KeySchedule_buffer3_amount(KeySchedule_buffer3_amount),
         .valid(memoryMappedEnable[6]),
         .wstrb(wstrb),
         .addr(addr[8:0]),
         .rdata(unitRData[6]),
         .ready(unitReady[6]),
         .wdata(wdata),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         KeySchedule  key7_17 (
         .out0(output_49_0),
         .out1(output_49_1),
         .out2(output_49_2),
         .out3(output_49_3),
         .out4(output_49_4),
         .out5(output_49_5),
         .out6(output_49_6),
         .out7(output_49_7),
         .out8(output_49_8),
         .out9(output_49_9),
         .out10(output_49_10),
         .out11(output_49_11),
         .out12(output_49_12),
         .out13(output_49_13),
         .out14(output_49_14),
         .out15(output_49_15),
         .in16(output_39_0),
         .in0(output_94_0),
         .in1(output_95_0),
         .in2(output_96_0),
         .in3(output_97_0),
         .in4(output_98_0),
         .in5(output_99_0),
         .in6(output_100_0),
         .in7(output_101_0),
         .in8(output_102_0),
         .in9(output_103_0),
         .in10(output_104_0),
         .in11(output_105_0),
         .in12(output_106_0),
         .in13(output_107_0),
         .in14(output_108_0),
         .in15(output_109_0),
         .KeySchedule_buffer0_amount(KeySchedule_buffer0_amount),
         .KeySchedule_buffer1_amount(KeySchedule_buffer1_amount),
         .KeySchedule_buffer2_amount(KeySchedule_buffer2_amount),
         .KeySchedule_buffer3_amount(KeySchedule_buffer3_amount),
         .valid(memoryMappedEnable[7]),
         .wstrb(wstrb),
         .addr(addr[8:0]),
         .rdata(unitRData[7]),
         .ready(unitReady[7]),
         .wdata(wdata),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         KeySchedule  key8_18 (
         .out0(output_50_0),
         .out1(output_50_1),
         .out2(output_50_2),
         .out3(output_50_3),
         .out4(output_50_4),
         .out5(output_50_5),
         .out6(output_50_6),
         .out7(output_50_7),
         .out8(output_50_8),
         .out9(output_50_9),
         .out10(output_50_10),
         .out11(output_50_11),
         .out12(output_50_12),
         .out13(output_50_13),
         .out14(output_50_14),
         .out15(output_50_15),
         .in16(output_40_0),
         .in0(output_78_0),
         .in1(output_79_0),
         .in2(output_80_0),
         .in3(output_81_0),
         .in4(output_82_0),
         .in5(output_83_0),
         .in6(output_84_0),
         .in7(output_85_0),
         .in8(output_86_0),
         .in9(output_87_0),
         .in10(output_88_0),
         .in11(output_89_0),
         .in12(output_90_0),
         .in13(output_91_0),
         .in14(output_92_0),
         .in15(output_93_0),
         .KeySchedule_buffer0_amount(KeySchedule_buffer0_amount),
         .KeySchedule_buffer1_amount(KeySchedule_buffer1_amount),
         .KeySchedule_buffer2_amount(KeySchedule_buffer2_amount),
         .KeySchedule_buffer3_amount(KeySchedule_buffer3_amount),
         .valid(memoryMappedEnable[8]),
         .wstrb(wstrb),
         .addr(addr[8:0]),
         .rdata(unitRData[8]),
         .ready(unitReady[8]),
         .wdata(wdata),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         KeySchedule  key9_19 (
         .out0(output_51_0),
         .out1(output_51_1),
         .out2(output_51_2),
         .out3(output_51_3),
         .out4(output_51_4),
         .out5(output_51_5),
         .out6(output_51_6),
         .out7(output_51_7),
         .out8(output_51_8),
         .out9(output_51_9),
         .out10(output_51_10),
         .out11(output_51_11),
         .out12(output_51_12),
         .out13(output_51_13),
         .out14(output_51_14),
         .out15(output_51_15),
         .in3(output_50_3),
         .in7(output_50_7),
         .in11(output_50_11),
         .in15(output_50_15),
         .in16(output_41_0),
         .in0(output_66_0),
         .in1(output_67_0),
         .in2(output_68_0),
         .in4(output_69_0),
         .in5(output_70_0),
         .in6(output_71_0),
         .in8(output_72_0),
         .in9(output_73_0),
         .in10(output_74_0),
         .in12(output_75_0),
         .in13(output_76_0),
         .in14(output_77_0),
         .KeySchedule_buffer0_amount(KeySchedule_buffer0_amount),
         .KeySchedule_buffer1_amount(KeySchedule_buffer1_amount),
         .KeySchedule_buffer2_amount(KeySchedule_buffer2_amount),
         .KeySchedule_buffer3_amount(KeySchedule_buffer3_amount),
         .valid(memoryMappedEnable[9]),
         .wstrb(wstrb),
         .addr(addr[8:0]),
         .rdata(unitRData[9]),
         .ready(unitReady[9]),
         .wdata(wdata),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         AddRoundKey  firstKey_20 (
         .out0(output_52_0),
         .out1(output_52_1),
         .out2(output_52_2),
         .out3(output_52_3),
         .out4(output_52_4),
         .out5(output_52_5),
         .out6(output_52_6),
         .out7(output_52_7),
         .out8(output_52_8),
         .out9(output_52_9),
         .out10(output_52_10),
         .out11(output_52_11),
         .out12(output_52_12),
         .out13(output_52_13),
         .out14(output_52_14),
         .out15(output_52_15),
         .in0(in0), // x0
         .in1(in1), // x1
         .in2(in2), // x2
         .in3(in3), // x3
         .in4(in4), // x4
         .in5(in5), // x5
         .in6(in6), // x6
         .in7(in7), // x7
         .in8(in8), // x8
         .in9(in9), // x9
         .in10(in10), // xa
         .in11(in11), // xb
         .in12(in12), // xc
         .in13(in13), // xd
         .in14(in14), // xe
         .in15(in15), // xf
         .in16(in16), // k0
         .in17(in17), // k1
         .in18(in18), // k2
         .in19(in19), // k3
         .in20(in20), // k4
         .in21(in21), // k5
         .in22(in22), // k6
         .in23(in23), // k7
         .in24(in24), // k8
         .in25(in25), // k9
         .in26(in26), // ka
         .in27(in27), // kb
         .in28(in28), // kc
         .in29(in29), // kd
         .in30(in30), // ke
         .in31(in31), // kf
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         MainRound  round0_21 (
         .out0(output_53_0),
         .out1(output_53_1),
         .out2(output_53_2),
         .out3(output_53_3),
         .out4(output_53_4),
         .out5(output_53_5),
         .out6(output_53_6),
         .out7(output_53_7),
         .out8(output_53_8),
         .out9(output_53_9),
         .out10(output_53_10),
         .out11(output_53_11),
         .out12(output_53_12),
         .out13(output_53_13),
         .out14(output_53_14),
         .out15(output_53_15),
         .in0(output_52_0),
         .in1(output_52_1),
         .in2(output_52_2),
         .in3(output_52_3),
         .in4(output_52_4),
         .in5(output_52_5),
         .in6(output_52_6),
         .in7(output_52_7),
         .in8(output_52_8),
         .in9(output_52_9),
         .in10(output_52_10),
         .in11(output_52_11),
         .in12(output_52_12),
         .in13(output_52_13),
         .in14(output_52_14),
         .in15(output_52_15),
         .in16(output_42_0),
         .in17(output_42_1),
         .in18(output_42_2),
         .in19(output_42_3),
         .in20(output_42_4),
         .in21(output_42_5),
         .in22(output_42_6),
         .in23(output_42_7),
         .in24(output_42_8),
         .in25(output_42_9),
         .in26(output_42_10),
         .in27(output_42_11),
         .in28(output_42_12),
         .in29(output_42_13),
         .in30(output_42_14),
         .in31(output_42_15),
         .DoRow_buffer0_amount(DoRow_buffer0_amount),
         .DoRow_buffer1_amount(DoRow_buffer1_amount),
         .DoRow_buffer2_amount(DoRow_buffer2_amount),
         .DoRow_buffer3_amount(DoRow_buffer3_amount),
         .DoRow_buffer4_amount(DoRow_buffer4_amount),
         .DoRow_buffer5_amount(DoRow_buffer5_amount),
         .DoRow_buffer6_amount(DoRow_buffer6_amount),
         .DoRow_buffer7_amount(DoRow_buffer7_amount),
         .valid(memoryMappedEnable[10]),
         .wstrb(wstrb),
         .addr(addr[12:0]),
         .rdata(unitRData[10]),
         .ready(unitReady[10]),
         .wdata(wdata),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         MainRound  round1_22 (
         .out0(output_54_0),
         .out1(output_54_1),
         .out2(output_54_2),
         .out3(output_54_3),
         .out4(output_54_4),
         .out5(output_54_5),
         .out6(output_54_6),
         .out7(output_54_7),
         .out8(output_54_8),
         .out9(output_54_9),
         .out10(output_54_10),
         .out11(output_54_11),
         .out12(output_54_12),
         .out13(output_54_13),
         .out14(output_54_14),
         .out15(output_54_15),
         .in0(output_53_0),
         .in1(output_53_1),
         .in2(output_53_2),
         .in3(output_53_3),
         .in4(output_53_4),
         .in5(output_53_5),
         .in6(output_53_6),
         .in7(output_53_7),
         .in8(output_53_8),
         .in9(output_53_9),
         .in10(output_53_10),
         .in11(output_53_11),
         .in12(output_53_12),
         .in13(output_53_13),
         .in14(output_53_14),
         .in15(output_53_15),
         .in16(output_43_0),
         .in17(output_43_1),
         .in18(output_43_2),
         .in19(output_43_3),
         .in20(output_43_4),
         .in21(output_43_5),
         .in22(output_43_6),
         .in23(output_43_7),
         .in24(output_43_8),
         .in25(output_43_9),
         .in26(output_43_10),
         .in27(output_43_11),
         .in28(output_43_12),
         .in29(output_43_13),
         .in30(output_43_14),
         .in31(output_43_15),
         .DoRow_buffer0_amount(DoRow_buffer0_amount),
         .DoRow_buffer1_amount(DoRow_buffer1_amount),
         .DoRow_buffer2_amount(DoRow_buffer2_amount),
         .DoRow_buffer3_amount(DoRow_buffer3_amount),
         .DoRow_buffer4_amount(DoRow_buffer4_amount),
         .DoRow_buffer5_amount(DoRow_buffer5_amount),
         .DoRow_buffer6_amount(DoRow_buffer6_amount),
         .DoRow_buffer7_amount(DoRow_buffer7_amount),
         .valid(memoryMappedEnable[11]),
         .wstrb(wstrb),
         .addr(addr[12:0]),
         .rdata(unitRData[11]),
         .ready(unitReady[11]),
         .wdata(wdata),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         MainRound  round2_23 (
         .out0(output_55_0),
         .out1(output_55_1),
         .out2(output_55_2),
         .out3(output_55_3),
         .out4(output_55_4),
         .out5(output_55_5),
         .out6(output_55_6),
         .out7(output_55_7),
         .out8(output_55_8),
         .out9(output_55_9),
         .out10(output_55_10),
         .out11(output_55_11),
         .out12(output_55_12),
         .out13(output_55_13),
         .out14(output_55_14),
         .out15(output_55_15),
         .in0(output_54_0),
         .in1(output_54_1),
         .in2(output_54_2),
         .in3(output_54_3),
         .in4(output_54_4),
         .in5(output_54_5),
         .in6(output_54_6),
         .in7(output_54_7),
         .in8(output_54_8),
         .in9(output_54_9),
         .in10(output_54_10),
         .in11(output_54_11),
         .in12(output_54_12),
         .in13(output_54_13),
         .in14(output_54_14),
         .in15(output_54_15),
         .in16(output_44_0),
         .in17(output_44_1),
         .in18(output_44_2),
         .in19(output_44_3),
         .in20(output_44_4),
         .in21(output_44_5),
         .in22(output_44_6),
         .in23(output_44_7),
         .in24(output_44_8),
         .in25(output_44_9),
         .in26(output_44_10),
         .in27(output_44_11),
         .in28(output_44_12),
         .in29(output_44_13),
         .in30(output_44_14),
         .in31(output_44_15),
         .DoRow_buffer0_amount(DoRow_buffer0_amount),
         .DoRow_buffer1_amount(DoRow_buffer1_amount),
         .DoRow_buffer2_amount(DoRow_buffer2_amount),
         .DoRow_buffer3_amount(DoRow_buffer3_amount),
         .DoRow_buffer4_amount(DoRow_buffer4_amount),
         .DoRow_buffer5_amount(DoRow_buffer5_amount),
         .DoRow_buffer6_amount(DoRow_buffer6_amount),
         .DoRow_buffer7_amount(DoRow_buffer7_amount),
         .valid(memoryMappedEnable[12]),
         .wstrb(wstrb),
         .addr(addr[12:0]),
         .rdata(unitRData[12]),
         .ready(unitReady[12]),
         .wdata(wdata),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         MainRound  round3_24 (
         .out0(output_56_0),
         .out1(output_56_1),
         .out2(output_56_2),
         .out3(output_56_3),
         .out4(output_56_4),
         .out5(output_56_5),
         .out6(output_56_6),
         .out7(output_56_7),
         .out8(output_56_8),
         .out9(output_56_9),
         .out10(output_56_10),
         .out11(output_56_11),
         .out12(output_56_12),
         .out13(output_56_13),
         .out14(output_56_14),
         .out15(output_56_15),
         .in0(output_55_0),
         .in1(output_55_1),
         .in2(output_55_2),
         .in3(output_55_3),
         .in4(output_55_4),
         .in5(output_55_5),
         .in6(output_55_6),
         .in7(output_55_7),
         .in8(output_55_8),
         .in9(output_55_9),
         .in10(output_55_10),
         .in11(output_55_11),
         .in12(output_55_12),
         .in13(output_55_13),
         .in14(output_55_14),
         .in15(output_55_15),
         .in16(output_45_0),
         .in17(output_45_1),
         .in18(output_45_2),
         .in19(output_45_3),
         .in20(output_45_4),
         .in21(output_45_5),
         .in22(output_45_6),
         .in23(output_45_7),
         .in24(output_45_8),
         .in25(output_45_9),
         .in26(output_45_10),
         .in27(output_45_11),
         .in28(output_45_12),
         .in29(output_45_13),
         .in30(output_45_14),
         .in31(output_45_15),
         .DoRow_buffer0_amount(DoRow_buffer0_amount),
         .DoRow_buffer1_amount(DoRow_buffer1_amount),
         .DoRow_buffer2_amount(DoRow_buffer2_amount),
         .DoRow_buffer3_amount(DoRow_buffer3_amount),
         .DoRow_buffer4_amount(DoRow_buffer4_amount),
         .DoRow_buffer5_amount(DoRow_buffer5_amount),
         .DoRow_buffer6_amount(DoRow_buffer6_amount),
         .DoRow_buffer7_amount(DoRow_buffer7_amount),
         .valid(memoryMappedEnable[13]),
         .wstrb(wstrb),
         .addr(addr[12:0]),
         .rdata(unitRData[13]),
         .ready(unitReady[13]),
         .wdata(wdata),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         MainRound  round4_25 (
         .out0(output_57_0),
         .out1(output_57_1),
         .out2(output_57_2),
         .out3(output_57_3),
         .out4(output_57_4),
         .out5(output_57_5),
         .out6(output_57_6),
         .out7(output_57_7),
         .out8(output_57_8),
         .out9(output_57_9),
         .out10(output_57_10),
         .out11(output_57_11),
         .out12(output_57_12),
         .out13(output_57_13),
         .out14(output_57_14),
         .out15(output_57_15),
         .in0(output_56_0),
         .in1(output_56_1),
         .in2(output_56_2),
         .in3(output_56_3),
         .in4(output_56_4),
         .in5(output_56_5),
         .in6(output_56_6),
         .in7(output_56_7),
         .in8(output_56_8),
         .in9(output_56_9),
         .in10(output_56_10),
         .in11(output_56_11),
         .in12(output_56_12),
         .in13(output_56_13),
         .in14(output_56_14),
         .in15(output_56_15),
         .in16(output_46_0),
         .in17(output_46_1),
         .in18(output_46_2),
         .in19(output_46_3),
         .in20(output_46_4),
         .in21(output_46_5),
         .in22(output_46_6),
         .in23(output_46_7),
         .in24(output_46_8),
         .in25(output_46_9),
         .in26(output_46_10),
         .in27(output_46_11),
         .in28(output_46_12),
         .in29(output_46_13),
         .in30(output_46_14),
         .in31(output_46_15),
         .DoRow_buffer0_amount(DoRow_buffer0_amount),
         .DoRow_buffer1_amount(DoRow_buffer1_amount),
         .DoRow_buffer2_amount(DoRow_buffer2_amount),
         .DoRow_buffer3_amount(DoRow_buffer3_amount),
         .DoRow_buffer4_amount(DoRow_buffer4_amount),
         .DoRow_buffer5_amount(DoRow_buffer5_amount),
         .DoRow_buffer6_amount(DoRow_buffer6_amount),
         .DoRow_buffer7_amount(DoRow_buffer7_amount),
         .valid(memoryMappedEnable[14]),
         .wstrb(wstrb),
         .addr(addr[12:0]),
         .rdata(unitRData[14]),
         .ready(unitReady[14]),
         .wdata(wdata),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         MainRound  round5_26 (
         .out0(output_58_0),
         .out1(output_58_1),
         .out2(output_58_2),
         .out3(output_58_3),
         .out4(output_58_4),
         .out5(output_58_5),
         .out6(output_58_6),
         .out7(output_58_7),
         .out8(output_58_8),
         .out9(output_58_9),
         .out10(output_58_10),
         .out11(output_58_11),
         .out12(output_58_12),
         .out13(output_58_13),
         .out14(output_58_14),
         .out15(output_58_15),
         .in0(output_57_0),
         .in1(output_57_1),
         .in2(output_57_2),
         .in3(output_57_3),
         .in4(output_57_4),
         .in5(output_57_5),
         .in6(output_57_6),
         .in7(output_57_7),
         .in8(output_57_8),
         .in9(output_57_9),
         .in10(output_57_10),
         .in11(output_57_11),
         .in12(output_57_12),
         .in13(output_57_13),
         .in14(output_57_14),
         .in15(output_57_15),
         .in16(output_47_0),
         .in17(output_47_1),
         .in18(output_47_2),
         .in19(output_47_3),
         .in20(output_47_4),
         .in21(output_47_5),
         .in22(output_47_6),
         .in23(output_47_7),
         .in24(output_47_8),
         .in25(output_47_9),
         .in26(output_47_10),
         .in27(output_47_11),
         .in28(output_47_12),
         .in29(output_47_13),
         .in30(output_47_14),
         .in31(output_47_15),
         .DoRow_buffer0_amount(DoRow_buffer0_amount),
         .DoRow_buffer1_amount(DoRow_buffer1_amount),
         .DoRow_buffer2_amount(DoRow_buffer2_amount),
         .DoRow_buffer3_amount(DoRow_buffer3_amount),
         .DoRow_buffer4_amount(DoRow_buffer4_amount),
         .DoRow_buffer5_amount(DoRow_buffer5_amount),
         .DoRow_buffer6_amount(DoRow_buffer6_amount),
         .DoRow_buffer7_amount(DoRow_buffer7_amount),
         .valid(memoryMappedEnable[15]),
         .wstrb(wstrb),
         .addr(addr[12:0]),
         .rdata(unitRData[15]),
         .ready(unitReady[15]),
         .wdata(wdata),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         MainRound  round6_27 (
         .out0(output_59_0),
         .out1(output_59_1),
         .out2(output_59_2),
         .out3(output_59_3),
         .out4(output_59_4),
         .out5(output_59_5),
         .out6(output_59_6),
         .out7(output_59_7),
         .out8(output_59_8),
         .out9(output_59_9),
         .out10(output_59_10),
         .out11(output_59_11),
         .out12(output_59_12),
         .out13(output_59_13),
         .out14(output_59_14),
         .out15(output_59_15),
         .in0(output_58_0),
         .in1(output_58_1),
         .in2(output_58_2),
         .in3(output_58_3),
         .in4(output_58_4),
         .in5(output_58_5),
         .in6(output_58_6),
         .in7(output_58_7),
         .in8(output_58_8),
         .in9(output_58_9),
         .in10(output_58_10),
         .in11(output_58_11),
         .in12(output_58_12),
         .in13(output_58_13),
         .in14(output_58_14),
         .in15(output_58_15),
         .in16(output_48_0),
         .in17(output_48_1),
         .in18(output_48_2),
         .in19(output_48_3),
         .in20(output_48_4),
         .in21(output_48_5),
         .in22(output_48_6),
         .in23(output_48_7),
         .in24(output_48_8),
         .in25(output_48_9),
         .in26(output_48_10),
         .in27(output_48_11),
         .in28(output_48_12),
         .in29(output_48_13),
         .in30(output_48_14),
         .in31(output_48_15),
         .DoRow_buffer0_amount(DoRow_buffer0_amount),
         .DoRow_buffer1_amount(DoRow_buffer1_amount),
         .DoRow_buffer2_amount(DoRow_buffer2_amount),
         .DoRow_buffer3_amount(DoRow_buffer3_amount),
         .DoRow_buffer4_amount(DoRow_buffer4_amount),
         .DoRow_buffer5_amount(DoRow_buffer5_amount),
         .DoRow_buffer6_amount(DoRow_buffer6_amount),
         .DoRow_buffer7_amount(DoRow_buffer7_amount),
         .valid(memoryMappedEnable[16]),
         .wstrb(wstrb),
         .addr(addr[12:0]),
         .rdata(unitRData[16]),
         .ready(unitReady[16]),
         .wdata(wdata),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         MainRound  round7_28 (
         .out0(output_60_0),
         .out1(output_60_1),
         .out2(output_60_2),
         .out3(output_60_3),
         .out4(output_60_4),
         .out5(output_60_5),
         .out6(output_60_6),
         .out7(output_60_7),
         .out8(output_60_8),
         .out9(output_60_9),
         .out10(output_60_10),
         .out11(output_60_11),
         .out12(output_60_12),
         .out13(output_60_13),
         .out14(output_60_14),
         .out15(output_60_15),
         .in0(output_59_0),
         .in1(output_59_1),
         .in2(output_59_2),
         .in3(output_59_3),
         .in4(output_59_4),
         .in5(output_59_5),
         .in6(output_59_6),
         .in7(output_59_7),
         .in8(output_59_8),
         .in9(output_59_9),
         .in10(output_59_10),
         .in11(output_59_11),
         .in12(output_59_12),
         .in13(output_59_13),
         .in14(output_59_14),
         .in15(output_59_15),
         .in16(output_49_0),
         .in17(output_49_1),
         .in18(output_49_2),
         .in19(output_49_3),
         .in20(output_49_4),
         .in21(output_49_5),
         .in22(output_49_6),
         .in23(output_49_7),
         .in24(output_49_8),
         .in25(output_49_9),
         .in26(output_49_10),
         .in27(output_49_11),
         .in28(output_49_12),
         .in29(output_49_13),
         .in30(output_49_14),
         .in31(output_49_15),
         .DoRow_buffer0_amount(DoRow_buffer0_amount),
         .DoRow_buffer1_amount(DoRow_buffer1_amount),
         .DoRow_buffer2_amount(DoRow_buffer2_amount),
         .DoRow_buffer3_amount(DoRow_buffer3_amount),
         .DoRow_buffer4_amount(DoRow_buffer4_amount),
         .DoRow_buffer5_amount(DoRow_buffer5_amount),
         .DoRow_buffer6_amount(DoRow_buffer6_amount),
         .DoRow_buffer7_amount(DoRow_buffer7_amount),
         .valid(memoryMappedEnable[17]),
         .wstrb(wstrb),
         .addr(addr[12:0]),
         .rdata(unitRData[17]),
         .ready(unitReady[17]),
         .wdata(wdata),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         MainRound  round8_29 (
         .out0(output_61_0),
         .out1(output_61_1),
         .out2(output_61_2),
         .out3(output_61_3),
         .out4(output_61_4),
         .out5(output_61_5),
         .out6(output_61_6),
         .out7(output_61_7),
         .out8(output_61_8),
         .out9(output_61_9),
         .out10(output_61_10),
         .out11(output_61_11),
         .out12(output_61_12),
         .out13(output_61_13),
         .out14(output_61_14),
         .out15(output_61_15),
         .in0(output_60_0),
         .in1(output_60_1),
         .in2(output_60_2),
         .in3(output_60_3),
         .in4(output_60_4),
         .in5(output_60_5),
         .in6(output_60_6),
         .in7(output_60_7),
         .in8(output_60_8),
         .in9(output_60_9),
         .in10(output_60_10),
         .in11(output_60_11),
         .in12(output_60_12),
         .in13(output_60_13),
         .in14(output_60_14),
         .in15(output_60_15),
         .in16(output_50_0),
         .in17(output_50_1),
         .in18(output_50_2),
         .in19(output_50_3),
         .in20(output_50_4),
         .in21(output_50_5),
         .in22(output_50_6),
         .in23(output_50_7),
         .in24(output_50_8),
         .in25(output_50_9),
         .in26(output_50_10),
         .in27(output_50_11),
         .in28(output_50_12),
         .in29(output_50_13),
         .in30(output_50_14),
         .in31(output_50_15),
         .DoRow_buffer0_amount(DoRow_buffer0_amount),
         .DoRow_buffer1_amount(DoRow_buffer1_amount),
         .DoRow_buffer2_amount(DoRow_buffer2_amount),
         .DoRow_buffer3_amount(DoRow_buffer3_amount),
         .DoRow_buffer4_amount(DoRow_buffer4_amount),
         .DoRow_buffer5_amount(DoRow_buffer5_amount),
         .DoRow_buffer6_amount(DoRow_buffer6_amount),
         .DoRow_buffer7_amount(DoRow_buffer7_amount),
         .valid(memoryMappedEnable[18]),
         .wstrb(wstrb),
         .addr(addr[12:0]),
         .rdata(unitRData[18]),
         .ready(unitReady[18]),
         .wdata(wdata),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         SBox  subBytes_30 (
         .out0(output_62_0),
         .out1(output_62_1),
         .out2(output_62_2),
         .out3(output_62_3),
         .out4(output_62_4),
         .out5(output_62_5),
         .out6(output_62_6),
         .out7(output_62_7),
         .out8(output_62_8),
         .out9(output_62_9),
         .out10(output_62_10),
         .out11(output_62_11),
         .out12(output_62_12),
         .out13(output_62_13),
         .out14(output_62_14),
         .out15(output_62_15),
         .in0(output_61_0),
         .in1(output_61_1),
         .in2(output_61_2),
         .in3(output_61_3),
         .in4(output_61_4),
         .in5(output_61_5),
         .in6(output_61_6),
         .in7(output_61_7),
         .in8(output_61_8),
         .in9(output_61_9),
         .in10(output_61_10),
         .in11(output_61_11),
         .in12(output_61_12),
         .in13(output_61_13),
         .in14(output_61_14),
         .in15(output_61_15),
         .valid(memoryMappedEnable[19]),
         .wstrb(wstrb),
         .addr(addr[10:0]),
         .rdata(unitRData[19]),
         .ready(unitReady[19]),
         .wdata(wdata),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         ShiftRows  shiftRows_31 (
         .out0(output_63_0),
         .out1(output_63_1),
         .out2(output_63_2),
         .out3(output_63_3),
         .out4(output_63_4),
         .out5(output_63_5),
         .out6(output_63_6),
         .out7(output_63_7),
         .out8(output_63_8),
         .out9(output_63_9),
         .out10(output_63_10),
         .out11(output_63_11),
         .out12(output_63_12),
         .out13(output_63_13),
         .out14(output_63_14),
         .out15(output_63_15),
         .in0(output_62_0),
         .in1(output_62_1),
         .in2(output_62_2),
         .in3(output_62_3),
         .in4(output_62_4),
         .in5(output_62_5),
         .in6(output_62_6),
         .in7(output_62_7),
         .in8(output_62_8),
         .in9(output_62_9),
         .in10(output_62_10),
         .in11(output_62_11),
         .in12(output_62_12),
         .in13(output_62_13),
         .in14(output_62_14),
         .in15(output_62_15),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         AddRoundKey  lastKey_32 (
         .out0(output_64_0),
         .out1(output_64_1),
         .out2(output_64_2),
         .out3(output_64_3),
         .out4(output_64_4),
         .out5(output_64_5),
         .out6(output_64_6),
         .out7(output_64_7),
         .out8(output_64_8),
         .out9(output_64_9),
         .out10(output_64_10),
         .out11(output_64_11),
         .out12(output_64_12),
         .out13(output_64_13),
         .out14(output_64_14),
         .out15(output_64_15),
         .in0(output_63_0),
         .in1(output_63_1),
         .in2(output_63_2),
         .in3(output_63_3),
         .in4(output_63_4),
         .in5(output_63_5),
         .in6(output_63_6),
         .in7(output_63_7),
         .in8(output_63_8),
         .in9(output_63_9),
         .in10(output_63_10),
         .in11(output_63_11),
         .in12(output_63_12),
         .in13(output_63_13),
         .in14(output_63_14),
         .in15(output_63_15),
         .in16(output_51_0),
         .in17(output_51_1),
         .in18(output_51_2),
         .in19(output_51_3),
         .in20(output_51_4),
         .in21(output_51_5),
         .in22(output_51_6),
         .in23(output_51_7),
         .in24(output_51_8),
         .in25(output_51_9),
         .in26(output_51_10),
         .in27(output_51_11),
         .in28(output_51_12),
         .in29(output_51_13),
         .in30(output_51_14),
         .in31(output_51_15),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer0_33 (
         .out0(output_66_0),
         .in0(output_50_0),
         .amount(AES_buffer0_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer1_34 (
         .out0(output_67_0),
         .in0(output_50_1),
         .amount(AES_buffer1_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer2_35 (
         .out0(output_68_0),
         .in0(output_50_2),
         .amount(AES_buffer2_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer3_36 (
         .out0(output_69_0),
         .in0(output_50_4),
         .amount(AES_buffer3_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer4_37 (
         .out0(output_70_0),
         .in0(output_50_5),
         .amount(AES_buffer4_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer5_38 (
         .out0(output_71_0),
         .in0(output_50_6),
         .amount(AES_buffer5_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer6_39 (
         .out0(output_72_0),
         .in0(output_50_8),
         .amount(AES_buffer6_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer7_40 (
         .out0(output_73_0),
         .in0(output_50_9),
         .amount(AES_buffer7_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer8_41 (
         .out0(output_74_0),
         .in0(output_50_10),
         .amount(AES_buffer8_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer9_42 (
         .out0(output_75_0),
         .in0(output_50_12),
         .amount(AES_buffer9_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer10_43 (
         .out0(output_76_0),
         .in0(output_50_13),
         .amount(AES_buffer10_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer11_44 (
         .out0(output_77_0),
         .in0(output_50_14),
         .amount(AES_buffer11_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer12_45 (
         .out0(output_78_0),
         .in0(output_49_0),
         .amount(AES_buffer12_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer13_46 (
         .out0(output_79_0),
         .in0(output_49_1),
         .amount(AES_buffer13_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer14_47 (
         .out0(output_80_0),
         .in0(output_49_2),
         .amount(AES_buffer14_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer15_48 (
         .out0(output_81_0),
         .in0(output_49_3),
         .amount(AES_buffer15_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer16_49 (
         .out0(output_82_0),
         .in0(output_49_4),
         .amount(AES_buffer16_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer17_50 (
         .out0(output_83_0),
         .in0(output_49_5),
         .amount(AES_buffer17_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer18_51 (
         .out0(output_84_0),
         .in0(output_49_6),
         .amount(AES_buffer18_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer19_52 (
         .out0(output_85_0),
         .in0(output_49_7),
         .amount(AES_buffer19_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer20_53 (
         .out0(output_86_0),
         .in0(output_49_8),
         .amount(AES_buffer20_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer21_54 (
         .out0(output_87_0),
         .in0(output_49_9),
         .amount(AES_buffer21_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer22_55 (
         .out0(output_88_0),
         .in0(output_49_10),
         .amount(AES_buffer22_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer23_56 (
         .out0(output_89_0),
         .in0(output_49_11),
         .amount(AES_buffer23_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer24_57 (
         .out0(output_90_0),
         .in0(output_49_12),
         .amount(AES_buffer24_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer25_58 (
         .out0(output_91_0),
         .in0(output_49_13),
         .amount(AES_buffer25_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer26_59 (
         .out0(output_92_0),
         .in0(output_49_14),
         .amount(AES_buffer26_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer27_60 (
         .out0(output_93_0),
         .in0(output_49_15),
         .amount(AES_buffer27_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer28_61 (
         .out0(output_94_0),
         .in0(output_48_0),
         .amount(AES_buffer28_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer29_62 (
         .out0(output_95_0),
         .in0(output_48_1),
         .amount(AES_buffer29_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer30_63 (
         .out0(output_96_0),
         .in0(output_48_2),
         .amount(AES_buffer30_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer31_64 (
         .out0(output_97_0),
         .in0(output_48_3),
         .amount(AES_buffer31_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer32_65 (
         .out0(output_98_0),
         .in0(output_48_4),
         .amount(AES_buffer32_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer33_66 (
         .out0(output_99_0),
         .in0(output_48_5),
         .amount(AES_buffer33_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer34_67 (
         .out0(output_100_0),
         .in0(output_48_6),
         .amount(AES_buffer34_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer35_68 (
         .out0(output_101_0),
         .in0(output_48_7),
         .amount(AES_buffer35_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer36_69 (
         .out0(output_102_0),
         .in0(output_48_8),
         .amount(AES_buffer36_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer37_70 (
         .out0(output_103_0),
         .in0(output_48_9),
         .amount(AES_buffer37_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer38_71 (
         .out0(output_104_0),
         .in0(output_48_10),
         .amount(AES_buffer38_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer39_72 (
         .out0(output_105_0),
         .in0(output_48_11),
         .amount(AES_buffer39_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer40_73 (
         .out0(output_106_0),
         .in0(output_48_12),
         .amount(AES_buffer40_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer41_74 (
         .out0(output_107_0),
         .in0(output_48_13),
         .amount(AES_buffer41_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer42_75 (
         .out0(output_108_0),
         .in0(output_48_14),
         .amount(AES_buffer42_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer43_76 (
         .out0(output_109_0),
         .in0(output_48_15),
         .amount(AES_buffer43_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer44_77 (
         .out0(output_110_0),
         .in0(output_47_0),
         .amount(AES_buffer44_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer45_78 (
         .out0(output_111_0),
         .in0(output_47_1),
         .amount(AES_buffer45_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer46_79 (
         .out0(output_112_0),
         .in0(output_47_2),
         .amount(AES_buffer46_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer47_80 (
         .out0(output_113_0),
         .in0(output_47_3),
         .amount(AES_buffer47_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer48_81 (
         .out0(output_114_0),
         .in0(output_47_4),
         .amount(AES_buffer48_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer49_82 (
         .out0(output_115_0),
         .in0(output_47_5),
         .amount(AES_buffer49_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer50_83 (
         .out0(output_116_0),
         .in0(output_47_6),
         .amount(AES_buffer50_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer51_84 (
         .out0(output_117_0),
         .in0(output_47_7),
         .amount(AES_buffer51_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer52_85 (
         .out0(output_118_0),
         .in0(output_47_8),
         .amount(AES_buffer52_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer53_86 (
         .out0(output_119_0),
         .in0(output_47_9),
         .amount(AES_buffer53_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer54_87 (
         .out0(output_120_0),
         .in0(output_47_10),
         .amount(AES_buffer54_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer55_88 (
         .out0(output_121_0),
         .in0(output_47_11),
         .amount(AES_buffer55_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer56_89 (
         .out0(output_122_0),
         .in0(output_47_12),
         .amount(AES_buffer56_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer57_90 (
         .out0(output_123_0),
         .in0(output_47_13),
         .amount(AES_buffer57_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer58_91 (
         .out0(output_124_0),
         .in0(output_47_14),
         .amount(AES_buffer58_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer59_92 (
         .out0(output_125_0),
         .in0(output_47_15),
         .amount(AES_buffer59_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer60_93 (
         .out0(output_126_0),
         .in0(output_46_0),
         .amount(AES_buffer60_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer61_94 (
         .out0(output_127_0),
         .in0(output_46_1),
         .amount(AES_buffer61_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer62_95 (
         .out0(output_128_0),
         .in0(output_46_2),
         .amount(AES_buffer62_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer63_96 (
         .out0(output_129_0),
         .in0(output_46_3),
         .amount(AES_buffer63_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer64_97 (
         .out0(output_130_0),
         .in0(output_46_4),
         .amount(AES_buffer64_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer65_98 (
         .out0(output_131_0),
         .in0(output_46_5),
         .amount(AES_buffer65_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer66_99 (
         .out0(output_132_0),
         .in0(output_46_6),
         .amount(AES_buffer66_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer67_100 (
         .out0(output_133_0),
         .in0(output_46_7),
         .amount(AES_buffer67_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer68_101 (
         .out0(output_134_0),
         .in0(output_46_8),
         .amount(AES_buffer68_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer69_102 (
         .out0(output_135_0),
         .in0(output_46_9),
         .amount(AES_buffer69_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer70_103 (
         .out0(output_136_0),
         .in0(output_46_10),
         .amount(AES_buffer70_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer71_104 (
         .out0(output_137_0),
         .in0(output_46_11),
         .amount(AES_buffer71_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer72_105 (
         .out0(output_138_0),
         .in0(output_46_12),
         .amount(AES_buffer72_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer73_106 (
         .out0(output_139_0),
         .in0(output_46_13),
         .amount(AES_buffer73_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer74_107 (
         .out0(output_140_0),
         .in0(output_46_14),
         .amount(AES_buffer74_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer75_108 (
         .out0(output_141_0),
         .in0(output_46_15),
         .amount(AES_buffer75_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer76_109 (
         .out0(output_142_0),
         .in0(output_45_0),
         .amount(AES_buffer76_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer77_110 (
         .out0(output_143_0),
         .in0(output_45_1),
         .amount(AES_buffer77_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer78_111 (
         .out0(output_144_0),
         .in0(output_45_2),
         .amount(AES_buffer78_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer79_112 (
         .out0(output_145_0),
         .in0(output_45_3),
         .amount(AES_buffer79_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer80_113 (
         .out0(output_146_0),
         .in0(output_45_4),
         .amount(AES_buffer80_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer81_114 (
         .out0(output_147_0),
         .in0(output_45_5),
         .amount(AES_buffer81_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer82_115 (
         .out0(output_148_0),
         .in0(output_45_6),
         .amount(AES_buffer82_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer83_116 (
         .out0(output_149_0),
         .in0(output_45_7),
         .amount(AES_buffer83_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer84_117 (
         .out0(output_150_0),
         .in0(output_45_8),
         .amount(AES_buffer84_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer85_118 (
         .out0(output_151_0),
         .in0(output_45_9),
         .amount(AES_buffer85_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer86_119 (
         .out0(output_152_0),
         .in0(output_45_10),
         .amount(AES_buffer86_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer87_120 (
         .out0(output_153_0),
         .in0(output_45_11),
         .amount(AES_buffer87_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer88_121 (
         .out0(output_154_0),
         .in0(output_45_12),
         .amount(AES_buffer88_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer89_122 (
         .out0(output_155_0),
         .in0(output_45_13),
         .amount(AES_buffer89_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer90_123 (
         .out0(output_156_0),
         .in0(output_45_14),
         .amount(AES_buffer90_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer91_124 (
         .out0(output_157_0),
         .in0(output_45_15),
         .amount(AES_buffer91_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer92_125 (
         .out0(output_158_0),
         .in0(output_44_0),
         .amount(AES_buffer92_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer93_126 (
         .out0(output_159_0),
         .in0(output_44_1),
         .amount(AES_buffer93_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer94_127 (
         .out0(output_160_0),
         .in0(output_44_2),
         .amount(AES_buffer94_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer95_128 (
         .out0(output_161_0),
         .in0(output_44_3),
         .amount(AES_buffer95_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer96_129 (
         .out0(output_162_0),
         .in0(output_44_4),
         .amount(AES_buffer96_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer97_130 (
         .out0(output_163_0),
         .in0(output_44_5),
         .amount(AES_buffer97_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer98_131 (
         .out0(output_164_0),
         .in0(output_44_6),
         .amount(AES_buffer98_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer99_132 (
         .out0(output_165_0),
         .in0(output_44_7),
         .amount(AES_buffer99_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer100_133 (
         .out0(output_166_0),
         .in0(output_44_8),
         .amount(AES_buffer100_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer101_134 (
         .out0(output_167_0),
         .in0(output_44_9),
         .amount(AES_buffer101_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer102_135 (
         .out0(output_168_0),
         .in0(output_44_10),
         .amount(AES_buffer102_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer103_136 (
         .out0(output_169_0),
         .in0(output_44_11),
         .amount(AES_buffer103_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer104_137 (
         .out0(output_170_0),
         .in0(output_44_12),
         .amount(AES_buffer104_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer105_138 (
         .out0(output_171_0),
         .in0(output_44_13),
         .amount(AES_buffer105_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer106_139 (
         .out0(output_172_0),
         .in0(output_44_14),
         .amount(AES_buffer106_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer107_140 (
         .out0(output_173_0),
         .in0(output_44_15),
         .amount(AES_buffer107_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer108_141 (
         .out0(output_174_0),
         .in0(output_43_0),
         .amount(AES_buffer108_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer109_142 (
         .out0(output_175_0),
         .in0(output_43_1),
         .amount(AES_buffer109_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer110_143 (
         .out0(output_176_0),
         .in0(output_43_2),
         .amount(AES_buffer110_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer111_144 (
         .out0(output_177_0),
         .in0(output_43_3),
         .amount(AES_buffer111_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer112_145 (
         .out0(output_178_0),
         .in0(output_43_4),
         .amount(AES_buffer112_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer113_146 (
         .out0(output_179_0),
         .in0(output_43_5),
         .amount(AES_buffer113_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer114_147 (
         .out0(output_180_0),
         .in0(output_43_6),
         .amount(AES_buffer114_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer115_148 (
         .out0(output_181_0),
         .in0(output_43_7),
         .amount(AES_buffer115_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer116_149 (
         .out0(output_182_0),
         .in0(output_43_8),
         .amount(AES_buffer116_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer117_150 (
         .out0(output_183_0),
         .in0(output_43_9),
         .amount(AES_buffer117_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer118_151 (
         .out0(output_184_0),
         .in0(output_43_10),
         .amount(AES_buffer118_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer119_152 (
         .out0(output_185_0),
         .in0(output_43_11),
         .amount(AES_buffer119_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer120_153 (
         .out0(output_186_0),
         .in0(output_43_12),
         .amount(AES_buffer120_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer121_154 (
         .out0(output_187_0),
         .in0(output_43_13),
         .amount(AES_buffer121_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer122_155 (
         .out0(output_188_0),
         .in0(output_43_14),
         .amount(AES_buffer122_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer123_156 (
         .out0(output_189_0),
         .in0(output_43_15),
         .amount(AES_buffer123_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer124_157 (
         .out0(output_190_0),
         .in0(output_42_0),
         .amount(AES_buffer124_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer125_158 (
         .out0(output_191_0),
         .in0(output_42_1),
         .amount(AES_buffer125_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer126_159 (
         .out0(output_192_0),
         .in0(output_42_2),
         .amount(AES_buffer126_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer127_160 (
         .out0(output_193_0),
         .in0(output_42_3),
         .amount(AES_buffer127_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer128_161 (
         .out0(output_194_0),
         .in0(output_42_4),
         .amount(AES_buffer128_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer129_162 (
         .out0(output_195_0),
         .in0(output_42_5),
         .amount(AES_buffer129_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer130_163 (
         .out0(output_196_0),
         .in0(output_42_6),
         .amount(AES_buffer130_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer131_164 (
         .out0(output_197_0),
         .in0(output_42_7),
         .amount(AES_buffer131_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer132_165 (
         .out0(output_198_0),
         .in0(output_42_8),
         .amount(AES_buffer132_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer133_166 (
         .out0(output_199_0),
         .in0(output_42_9),
         .amount(AES_buffer133_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer134_167 (
         .out0(output_200_0),
         .in0(output_42_10),
         .amount(AES_buffer134_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer135_168 (
         .out0(output_201_0),
         .in0(output_42_11),
         .amount(AES_buffer135_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer136_169 (
         .out0(output_202_0),
         .in0(output_42_12),
         .amount(AES_buffer136_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer137_170 (
         .out0(output_203_0),
         .in0(output_42_13),
         .amount(AES_buffer137_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer138_171 (
         .out0(output_204_0),
         .in0(output_42_14),
         .amount(AES_buffer138_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer139_172 (
         .out0(output_205_0),
         .in0(output_42_15),
         .amount(AES_buffer139_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer140_173 (
         .out0(output_206_0),
         .in0(in31), // kf
         .amount(AES_buffer140_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer141_174 (
         .out0(output_207_0),
         .in0(in30), // ke
         .amount(AES_buffer141_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer142_175 (
         .out0(output_208_0),
         .in0(in29), // kd
         .amount(AES_buffer142_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer143_176 (
         .out0(output_209_0),
         .in0(in28), // kc
         .amount(AES_buffer143_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer144_177 (
         .out0(output_210_0),
         .in0(in27), // kb
         .amount(AES_buffer144_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer145_178 (
         .out0(output_211_0),
         .in0(in26), // ka
         .amount(AES_buffer145_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer146_179 (
         .out0(output_212_0),
         .in0(in25), // k9
         .amount(AES_buffer146_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer147_180 (
         .out0(output_213_0),
         .in0(in24), // k8
         .amount(AES_buffer147_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer148_181 (
         .out0(output_214_0),
         .in0(in23), // k7
         .amount(AES_buffer148_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer149_182 (
         .out0(output_215_0),
         .in0(in22), // k6
         .amount(AES_buffer149_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer150_183 (
         .out0(output_216_0),
         .in0(in21), // k5
         .amount(AES_buffer150_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer151_184 (
         .out0(output_217_0),
         .in0(in20), // k4
         .amount(AES_buffer151_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer152_185 (
         .out0(output_218_0),
         .in0(in19), // k3
         .amount(AES_buffer152_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer153_186 (
         .out0(output_219_0),
         .in0(in18), // k2
         .amount(AES_buffer153_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer154_187 (
         .out0(output_220_0),
         .in0(in17), // k1
         .amount(AES_buffer154_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         Buffer  buffer155_188 (
         .out0(output_221_0),
         .in0(in16), // k0
         .amount(AES_buffer155_amount),
         .run(run),

         .clk(clk),
         .rst(rst)
      );
         assign out0 = output_64_0;
   assign out1 = output_64_1;
   assign out2 = output_64_2;
   assign out3 = output_64_3;
   assign out4 = output_64_4;
   assign out5 = output_64_5;
   assign out6 = output_64_6;
   assign out7 = output_64_7;
   assign out8 = output_64_8;
   assign out9 = output_64_9;
   assign out10 = output_64_10;
   assign out11 = output_64_11;
   assign out12 = output_64_12;
   assign out13 = output_64_13;
   assign out14 = output_64_14;
   assign out15 = output_64_15;
   endmodule
