	always @(posedge clk) begin
		case (addr)
			DATA_W'd0: r_data <= DATA_W'h00001137;
			DATA_W'd1: r_data <= DATA_W'h00010113;
			DATA_W'd2: r_data <= DATA_W'h446000ef;
			DATA_W'd3: r_data <= DATA_W'h0b374a89;
			DATA_W'd4: r_data <= DATA_W'h20232000;
			DATA_W'd5: r_data <= DATA_W'h9002015b;
			DATA_W'd6: r_data <= DATA_W'h97b34785;
			DATA_W'd7: r_data <= DATA_W'h97aa00b7;
			DATA_W'd8: r_data <= DATA_W'h28f02023;
			DATA_W'd9: r_data <= DATA_W'h27838082;
			DATA_W'd10: r_data <= DATA_W'h57882800;
			DATA_W'd11: r_data <= DATA_W'h27838082;
			DATA_W'd12: r_data <= DATA_W'h43c82800;
			DATA_W'd13: r_data <= DATA_W'h27838082;
			DATA_W'd14: r_data <= DATA_W'h47882800;
			DATA_W'd15: r_data <= DATA_W'h27838082;
			DATA_W'd16: r_data <= DATA_W'h47c82800;
			DATA_W'd17: r_data <= DATA_W'h27838082;
			DATA_W'd18: r_data <= DATA_W'h4b882800;
			DATA_W'd19: r_data <= DATA_W'h27838082;
			DATA_W'd20: r_data <= DATA_W'h4bc82800;
			DATA_W'd21: r_data <= DATA_W'h27838082;
			DATA_W'd22: r_data <= DATA_W'h4f882800;
			DATA_W'd23: r_data <= DATA_W'h27838082;
			DATA_W'd24: r_data <= DATA_W'h4fc82800;
			DATA_W'd25: r_data <= DATA_W'h27838082;
			DATA_W'd26: r_data <= DATA_W'h53882800;
			DATA_W'd27: r_data <= DATA_W'h27838082;
			DATA_W'd28: r_data <= DATA_W'h53c82800;
			DATA_W'd29: r_data <= DATA_W'h11418082;
			DATA_W'd30: r_data <= DATA_W'h22d1c606;
			DATA_W'd31: r_data <= DATA_W'h40b2dd7d;
			DATA_W'd32: r_data <= DATA_W'h80820141;
			DATA_W'd33: r_data <= DATA_W'hc4221141;
			DATA_W'd34: r_data <= DATA_W'h842ac606;
			DATA_W'd35: r_data <= DATA_W'hdd7d2a4d;
			DATA_W'd36: r_data <= DATA_W'h44228522;
			DATA_W'd37: r_data <= DATA_W'h014140b2;
			DATA_W'd38: r_data <= DATA_W'h1141a261;
			DATA_W'd39: r_data <= DATA_W'h2a55c606;
			DATA_W'd40: r_data <= DATA_W'h40b2dd7d;
			DATA_W'd41: r_data <= DATA_W'h80820141;
			DATA_W'd42: r_data <= DATA_W'hc6061141;
			DATA_W'd43: r_data <= DATA_W'hdd7d225d;
			DATA_W'd44: r_data <= DATA_W'h014140b2;
			DATA_W'd45: r_data <= DATA_W'h1141aa51;
			DATA_W'd46: r_data <= DATA_W'hc422c606;
			DATA_W'd47: r_data <= DATA_W'h22a1842e;
			DATA_W'd48: r_data <= DATA_W'h22a94505;
			DATA_W'd49: r_data <= DATA_W'h22994501;
			DATA_W'd50: r_data <= DATA_W'h22b18522;
			DATA_W'd51: r_data <= DATA_W'h2ab14505;
			DATA_W'd52: r_data <= DATA_W'h40b24422;
			DATA_W'd53: r_data <= DATA_W'h01414505;
			DATA_W'd54: r_data <= DATA_W'h1141aab1;
			DATA_W'd55: r_data <= DATA_W'hc6064511;
			DATA_W'd56: r_data <= DATA_W'h40b23755;
			DATA_W'd57: r_data <= DATA_W'hbf410141;
			DATA_W'd58: r_data <= DATA_W'hc4221141;
			DATA_W'd59: r_data <= DATA_W'h842ac606;
			DATA_W'd60: r_data <= DATA_W'h00044503;
			DATA_W'd61: r_data <= DATA_W'h40b2e509;
			DATA_W'd62: r_data <= DATA_W'h01414422;
			DATA_W'd63: r_data <= DATA_W'h04058082;
			DATA_W'd64: r_data <= DATA_W'hb7fd3751;
			DATA_W'd65: r_data <= DATA_W'hc4221141;
			DATA_W'd66: r_data <= DATA_W'h842ac606;
			DATA_W'd67: r_data <= DATA_W'h00044503;
			DATA_W'd68: r_data <= DATA_W'h3f8d0405;
			DATA_W'd69: r_data <= DATA_W'hfff44783;
			DATA_W'd70: r_data <= DATA_W'h40b2fbf5;
			DATA_W'd71: r_data <= DATA_W'h01414422;
			DATA_W'd72: r_data <= DATA_W'h11018082;
			DATA_W'd73: r_data <= DATA_W'hcc22c64e;
			DATA_W'd74: r_data <= DATA_W'h0513842a;
			DATA_W'd75: r_data <= DATA_W'hce062c80;
			DATA_W'd76: r_data <= DATA_W'hc84aca26;
			DATA_W'd77: r_data <= DATA_W'h3f4d892e;
			DATA_W'd78: r_data <= DATA_W'h2d400513;
			DATA_W'd79: r_data <= DATA_W'h45213775;
			DATA_W'd80: r_data <= DATA_W'h85223791;
			DATA_W'd81: r_data <= DATA_W'h378d37c1;
			DATA_W'd82: r_data <= DATA_W'h3fb984aa;
			DATA_W'd83: r_data <= DATA_W'h3fa9842a;
			DATA_W'd84: r_data <= DATA_W'h04220542;
			DATA_W'd85: r_data <= DATA_W'h3f898c49;
			DATA_W'd86: r_data <= DATA_W'h14938c45;
			DATA_W'd87: r_data <= DATA_W'h45190185;
			DATA_W'd88: r_data <= DATA_W'h370d8cc1;
			DATA_W'd89: r_data <= DATA_W'h10634401;
			DATA_W'd90: r_data <= DATA_W'h05130294;
			DATA_W'd91: r_data <= DATA_W'h3fad2c80;
			DATA_W'd92: r_data <= DATA_W'h2f400513;
			DATA_W'd93: r_data <= DATA_W'h40f23f95;
			DATA_W'd94: r_data <= DATA_W'h44628522;
			DATA_W'd95: r_data <= DATA_W'h494244d2;
			DATA_W'd96: r_data <= DATA_W'h610549b2;
			DATA_W'd97: r_data <= DATA_W'h370d8082;
			DATA_W'd98: r_data <= DATA_W'h008907b3;
			DATA_W'd99: r_data <= DATA_W'h00a78023;
			DATA_W'd100: r_data <= DATA_W'hbfd10405;
			DATA_W'd101: r_data <= DATA_W'hc64e1101;
			DATA_W'd102: r_data <= DATA_W'h84aaca26;
			DATA_W'd103: r_data <= DATA_W'h2c800513;
			DATA_W'd104: r_data <= DATA_W'hcc22ce06;
			DATA_W'd105: r_data <= DATA_W'h842ec84a;
			DATA_W'd106: r_data <= DATA_W'h3f3d8932;
			DATA_W'd107: r_data <= DATA_W'h30800513;
			DATA_W'd108: r_data <= DATA_W'h451d3f25;
			DATA_W'd109: r_data <= DATA_W'h85263dc1;
			DATA_W'd110: r_data <= DATA_W'h751337b1;
			DATA_W'd111: r_data <= DATA_W'h35d90ff4;
			DATA_W'd112: r_data <= DATA_W'h40845513;
			DATA_W'd113: r_data <= DATA_W'h0ff57513;
			DATA_W'd114: r_data <= DATA_W'h55133d75;
			DATA_W'd115: r_data <= DATA_W'h75134104;
			DATA_W'd116: r_data <= DATA_W'h3d4d0ff5;
			DATA_W'd117: r_data <= DATA_W'h01845513;
			DATA_W'd118: r_data <= DATA_W'h44813575;
			DATA_W'd119: r_data <= DATA_W'h0084ce63;
			DATA_W'd120: r_data <= DATA_W'h2c800513;
			DATA_W'd121: r_data <= DATA_W'h44623711;
			DATA_W'd122: r_data <= DATA_W'h44d240f2;
			DATA_W'd123: r_data <= DATA_W'h49b24942;
			DATA_W'd124: r_data <= DATA_W'h32400513;
			DATA_W'd125: r_data <= DATA_W'hbdcd6105;
			DATA_W'd126: r_data <= DATA_W'h009907b3;
			DATA_W'd127: r_data <= DATA_W'h0007c503;
			DATA_W'd128: r_data <= DATA_W'h35490485;
			DATA_W'd129: r_data <= DATA_W'h2c23bfe1;
			DATA_W'd130: r_data <= DATA_W'h808234a0;
			DATA_W'd131: r_data <= DATA_W'h35802783;
			DATA_W'd132: r_data <= DATA_W'h00a78023;
			DATA_W'd133: r_data <= DATA_W'h27838082;
			DATA_W'd134: r_data <= DATA_W'h91233580;
			DATA_W'd135: r_data <= DATA_W'h808200a7;
			DATA_W'd136: r_data <= DATA_W'h35802783;
			DATA_W'd137: r_data <= DATA_W'h00a78223;
			DATA_W'd138: r_data <= DATA_W'h27838082;
			DATA_W'd139: r_data <= DATA_W'h82a33580;
			DATA_W'd140: r_data <= DATA_W'h808200a7;
			DATA_W'd141: r_data <= DATA_W'h35802783;
			DATA_W'd142: r_data <= DATA_W'h00a78323;
			DATA_W'd143: r_data <= DATA_W'h27838082;
			DATA_W'd144: r_data <= DATA_W'hc5033580;
			DATA_W'd145: r_data <= DATA_W'h80820007;
			DATA_W'd146: r_data <= DATA_W'h35802783;
			DATA_W'd147: r_data <= DATA_W'h0047c503;
			DATA_W'd148: r_data <= DATA_W'h27838082;
			DATA_W'd149: r_data <= DATA_W'hc5033580;
			DATA_W'd150: r_data <= DATA_W'h80820017;
			DATA_W'd151: r_data <= DATA_W'h00050313;
			DATA_W'd152: r_data <= DATA_W'h00060e63;
			DATA_W'd153: r_data <= DATA_W'h00058383;
			DATA_W'd154: r_data <= DATA_W'h00730023;
			DATA_W'd155: r_data <= DATA_W'hfff60613;
			DATA_W'd156: r_data <= DATA_W'h00130313;
			DATA_W'd157: r_data <= DATA_W'h00158593;
			DATA_W'd158: r_data <= DATA_W'hfe0616e3;
			DATA_W'd159: r_data <= DATA_W'h00008067;
			DATA_W'd160: r_data <= DATA_W'h00000000;
			DATA_W'd161: r_data <= DATA_W'h3a434347;
			DATA_W'd162: r_data <= DATA_W'h35672820;
			DATA_W'd163: r_data <= DATA_W'h62343639;
			DATA_W'd164: r_data <= DATA_W'h37646335;
			DATA_W'd165: r_data <= DATA_W'h20293732;
			DATA_W'd166: r_data <= DATA_W'h312e3131;
			DATA_W'd167: r_data <= DATA_W'h4100302e;
			DATA_W'd168: r_data <= DATA_W'h00000025;
			DATA_W'd169: r_data <= DATA_W'h63736972;
			DATA_W'd170: r_data <= DATA_W'h1b010076;
			DATA_W'd171: r_data <= DATA_W'h04000000;
			DATA_W'd172: r_data <= DATA_W'h76720510;
			DATA_W'd173: r_data <= DATA_W'h32693233;
			DATA_W'd174: r_data <= DATA_W'h6d5f3070;
			DATA_W'd175: r_data <= DATA_W'h5f307032;
			DATA_W'd176: r_data <= DATA_W'h30703263;
			DATA_W'd177: r_data <= DATA_W'h00000000;
			DATA_W'd178: r_data <= DATA_W'h2d624f49;
			DATA_W'd179: r_data <= DATA_W'h54524155;
			DATA_W'd180: r_data <= DATA_W'h00000000;
			DATA_W'd181: r_data <= DATA_W'h6572203a;
			DATA_W'd182: r_data <= DATA_W'h73657571;
			DATA_W'd183: r_data <= DATA_W'h676e6974;
			DATA_W'd184: r_data <= DATA_W'h206f7420;
			DATA_W'd185: r_data <= DATA_W'h65636572;
			DATA_W'd186: r_data <= DATA_W'h20657669;
			DATA_W'd187: r_data <= DATA_W'h656c6966;
			DATA_W'd188: r_data <= DATA_W'h0000000a;
			DATA_W'd189: r_data <= DATA_W'h6966203a;
			DATA_W'd190: r_data <= DATA_W'h7220656c;
			DATA_W'd191: r_data <= DATA_W'h69656365;
			DATA_W'd192: r_data <= DATA_W'h0a646576;
			DATA_W'd193: r_data <= DATA_W'h00000000;
			DATA_W'd194: r_data <= DATA_W'h6572203a;
			DATA_W'd195: r_data <= DATA_W'h73657571;
			DATA_W'd196: r_data <= DATA_W'h676e6974;
			DATA_W'd197: r_data <= DATA_W'h206f7420;
			DATA_W'd198: r_data <= DATA_W'h646e6573;
			DATA_W'd199: r_data <= DATA_W'h6c696620;
			DATA_W'd200: r_data <= DATA_W'h00000a65;
			DATA_W'd201: r_data <= DATA_W'h6966203a;
			DATA_W'd202: r_data <= DATA_W'h7320656c;
			DATA_W'd203: r_data <= DATA_W'h0a746e65;
			DATA_W'd204: r_data <= DATA_W'h00254100;
			DATA_W'd205: r_data <= DATA_W'h69720000;
			DATA_W'd206: r_data <= DATA_W'h00766373;
			DATA_W'd207: r_data <= DATA_W'h00001b01;
			DATA_W'd208: r_data <= DATA_W'h05100400;
			DATA_W'd209: r_data <= DATA_W'h32337672;
			DATA_W'd210: r_data <= DATA_W'h30703269;
			DATA_W'd211: r_data <= DATA_W'h70326d5f;
			DATA_W'd212: r_data <= DATA_W'h32635f30;
			DATA_W'd213: r_data <= DATA_W'h00003070;
			DATA_W'd214: r_data <= DATA_W'h00000000;
			DATA_W'd215: r_data <= DATA_W'h00002541;
			DATA_W'd216: r_data <= DATA_W'h73697200;
			DATA_W'd217: r_data <= DATA_W'h01007663;
			DATA_W'd218: r_data <= DATA_W'h0000001b;
			DATA_W'd219: r_data <= DATA_W'h72051004;
			DATA_W'd220: r_data <= DATA_W'h69323376;
			DATA_W'd221: r_data <= DATA_W'h5f307032;
			DATA_W'd222: r_data <= DATA_W'h3070326d;
			DATA_W'd223: r_data <= DATA_W'h7032635f;
			DATA_W'd224: r_data <= DATA_W'h23410030;
			DATA_W'd225: r_data <= DATA_W'h72000000;
			DATA_W'd226: r_data <= DATA_W'h76637369;
			DATA_W'd227: r_data <= DATA_W'h00190100;
			DATA_W'd228: r_data <= DATA_W'h72050000;
			DATA_W'd229: r_data <= DATA_W'h69323376;
			DATA_W'd230: r_data <= DATA_W'h5f307032;
			DATA_W'd231: r_data <= DATA_W'h3070326d;
			DATA_W'd232: r_data <= DATA_W'h7032635f;
			DATA_W'd233: r_data <= DATA_W'h00000030;
			DATA_W'd234: r_data <= DATA_W'h2d624f49;
			DATA_W'd235: r_data <= DATA_W'h746f6f42;
			DATA_W'd236: r_data <= DATA_W'h64616f6c;
			DATA_W'd237: r_data <= DATA_W'h00007265;
			DATA_W'd238: r_data <= DATA_W'h6f63203a;
			DATA_W'd239: r_data <= DATA_W'h63656e6e;
			DATA_W'd240: r_data <= DATA_W'h21646574;
			DATA_W'd241: r_data <= DATA_W'h0000000a;
			DATA_W'd242: r_data <= DATA_W'h4444203a;
			DATA_W'd243: r_data <= DATA_W'h6e692052;
			DATA_W'd244: r_data <= DATA_W'h65737520;
			DATA_W'd245: r_data <= DATA_W'h0000000a;
			DATA_W'd246: r_data <= DATA_W'h7270203a;
			DATA_W'd247: r_data <= DATA_W'h6172676f;
			DATA_W'd248: r_data <= DATA_W'h6f74206d;
			DATA_W'd249: r_data <= DATA_W'h6e757220;
			DATA_W'd250: r_data <= DATA_W'h6f726620;
			DATA_W'd251: r_data <= DATA_W'h4444206d;
			DATA_W'd252: r_data <= DATA_W'h00000a52;
			DATA_W'd253: r_data <= DATA_W'h6f4c203a;
			DATA_W'd254: r_data <= DATA_W'h6e696461;
			DATA_W'd255: r_data <= DATA_W'h69662067;
			DATA_W'd256: r_data <= DATA_W'h61776d72;
			DATA_W'd257: r_data <= DATA_W'h2e2e6572;
			DATA_W'd258: r_data <= DATA_W'h00000a2e;
			DATA_W'd259: r_data <= DATA_W'h6552203a;
			DATA_W'd260: r_data <= DATA_W'h72617473;
			DATA_W'd261: r_data <= DATA_W'h50432074;
			DATA_W'd262: r_data <= DATA_W'h6f742055;
			DATA_W'd263: r_data <= DATA_W'h6e757220;
			DATA_W'd264: r_data <= DATA_W'h65737520;
			DATA_W'd265: r_data <= DATA_W'h72702072;
			DATA_W'd266: r_data <= DATA_W'h6172676f;
			DATA_W'd267: r_data <= DATA_W'h2e2e2e6d;
			DATA_W'd268: r_data <= DATA_W'h0000000a;
			DATA_W'd269: r_data <= DATA_W'h6d726966;
			DATA_W'd270: r_data <= DATA_W'h65726177;
			DATA_W'd271: r_data <= DATA_W'h6e69622e;
			DATA_W'd272: r_data <= DATA_W'h00000000;
			DATA_W'd273: r_data <= DATA_W'h77665f73;
			DATA_W'd274: r_data <= DATA_W'h6e69622e;
			DATA_W'd275: r_data <= DATA_W'h71790000;
			DATA_W'd276: r_data <= DATA_W'h053745d1;
			DATA_W'd277: r_data <= DATA_W'hd6064000;
			DATA_W'd278: r_data <= DATA_W'hd226d422;
			DATA_W'd279: r_data <= DATA_W'h33c539a9;
			DATA_W'd280: r_data <= DATA_W'h4515c119;
			DATA_W'd281: r_data <= DATA_W'h33f53105;
			DATA_W'd282: r_data <= DATA_W'h0513d97d;
			DATA_W'd283: r_data <= DATA_W'h39ad3a80;
			DATA_W'd284: r_data <= DATA_W'h3b800513;
			DATA_W'd285: r_data <= DATA_W'h05133995;
			DATA_W'd286: r_data <= DATA_W'h31bd3a80;
			DATA_W'd287: r_data <= DATA_W'h3c800513;
			DATA_W'd288: r_data <= DATA_W'h051331a5;
			DATA_W'd289: r_data <= DATA_W'h318d3a80;
			DATA_W'd290: r_data <= DATA_W'h3d800513;
			DATA_W'd291: r_data <= DATA_W'h463539b1;
			DATA_W'd292: r_data <= DATA_W'h43400593;
			DATA_W'd293: r_data <= DATA_W'h33d90808;
			DATA_W'd294: r_data <= DATA_W'h47a13901;
			DATA_W'd295: r_data <= DATA_W'h1d634481;
			DATA_W'd296: r_data <= DATA_W'h05b700f5;
			DATA_W'd297: r_data <= DATA_W'h08088000;
			DATA_W'd298: r_data <= DATA_W'h84aa39ad;
			DATA_W'd299: r_data <= DATA_W'h3a800513;
			DATA_W'd300: r_data <= DATA_W'h05133925;
			DATA_W'd301: r_data <= DATA_W'h390d3f40;
			DATA_W'd302: r_data <= DATA_W'h05934625;
			DATA_W'd303: r_data <= DATA_W'h00484440;
			DATA_W'd304: r_data <= DATA_W'hc4913b71;
			DATA_W'd305: r_data <= DATA_W'h80000637;
			DATA_W'd306: r_data <= DATA_W'h004885a6;
			DATA_W'd307: r_data <= DATA_W'h051331e1;
			DATA_W'd308: r_data <= DATA_W'h39193a80;
			DATA_W'd309: r_data <= DATA_W'h40c00513;
			DATA_W'd310: r_data <= DATA_W'h3e713901;
			DATA_W'd311: r_data <= DATA_W'hdd7d3e89;
			DATA_W'd312: r_data <= DATA_W'h542250b2;
			DATA_W'd313: r_data <= DATA_W'h45015492;
			DATA_W'd314: r_data <= DATA_W'h80826145;
			DATA_W'd315: r_data <= DATA_W'h00002541;
			DATA_W'd316: r_data <= DATA_W'h73697200;
			DATA_W'd317: r_data <= DATA_W'h01007663;
			DATA_W'd318: r_data <= DATA_W'h0000001b;
			DATA_W'd319: r_data <= DATA_W'h72051004;
			DATA_W'd320: r_data <= DATA_W'h69323376;
			DATA_W'd321: r_data <= DATA_W'h5f307032;
			DATA_W'd322: r_data <= DATA_W'h3070326d;
			DATA_W'd323: r_data <= DATA_W'h7032635f;
			DATA_W'd324: r_data <= DATA_W'h1e410030;
			DATA_W'd325: r_data <= DATA_W'h72000000;
			DATA_W'd326: r_data <= DATA_W'h76637369;
			DATA_W'd327: r_data <= DATA_W'h00140100;
			DATA_W'd328: r_data <= DATA_W'h72050000;
			DATA_W'd329: r_data <= DATA_W'h69323376;
			DATA_W'd330: r_data <= DATA_W'h5f307032;
			DATA_W'd331: r_data <= DATA_W'h3070326d;
			DATA_W'd332: r_data <= DATA_W'h00000000;
			DATA_W'd333: r_data <= DATA_W'h00000000;
			DATA_W'd334: r_data <= DATA_W'h00000000;
			DATA_W'd335: r_data <= DATA_W'h00000000;
			DATA_W'd336: r_data <= DATA_W'h00000000;
			DATA_W'd337: r_data <= DATA_W'h00000000;
			DATA_W'd338: r_data <= DATA_W'h00000000;
			DATA_W'd339: r_data <= DATA_W'h00000000;
			DATA_W'd340: r_data <= DATA_W'h00000000;
			DATA_W'd341: r_data <= DATA_W'h00000000;
			DATA_W'd342: r_data <= DATA_W'h00000000;
			DATA_W'd343: r_data <= DATA_W'h00000000;
			DATA_W'd344: r_data <= DATA_W'h00000000;
			DATA_W'd345: r_data <= DATA_W'h00000000;
			DATA_W'd346: r_data <= DATA_W'h00000000;
			DATA_W'd347: r_data <= DATA_W'h00000000;
			DATA_W'd348: r_data <= DATA_W'h00000000;
			DATA_W'd349: r_data <= DATA_W'h00000000;
			DATA_W'd350: r_data <= DATA_W'h00000000;
			DATA_W'd351: r_data <= DATA_W'h00000000;
			DATA_W'd352: r_data <= DATA_W'h00000000;
			DATA_W'd353: r_data <= DATA_W'h00000000;
			DATA_W'd354: r_data <= DATA_W'h00000000;
			DATA_W'd355: r_data <= DATA_W'h00000000;
			DATA_W'd356: r_data <= DATA_W'h00000000;
			DATA_W'd357: r_data <= DATA_W'h00000000;
			DATA_W'd358: r_data <= DATA_W'h00000000;
			DATA_W'd359: r_data <= DATA_W'h00000000;
			DATA_W'd360: r_data <= DATA_W'h00000000;
			DATA_W'd361: r_data <= DATA_W'h00000000;
			DATA_W'd362: r_data <= DATA_W'h00000000;
			DATA_W'd363: r_data <= DATA_W'h00000000;
			DATA_W'd364: r_data <= DATA_W'h00000000;
			DATA_W'd365: r_data <= DATA_W'h00000000;
			DATA_W'd366: r_data <= DATA_W'h00000000;
			DATA_W'd367: r_data <= DATA_W'h00000000;
			DATA_W'd368: r_data <= DATA_W'h00000000;
			DATA_W'd369: r_data <= DATA_W'h00000000;
			DATA_W'd370: r_data <= DATA_W'h00000000;
			DATA_W'd371: r_data <= DATA_W'h00000000;
			DATA_W'd372: r_data <= DATA_W'h00000000;
			DATA_W'd373: r_data <= DATA_W'h00000000;
			DATA_W'd374: r_data <= DATA_W'h00000000;
			DATA_W'd375: r_data <= DATA_W'h00000000;
			DATA_W'd376: r_data <= DATA_W'h00000000;
			DATA_W'd377: r_data <= DATA_W'h00000000;
			DATA_W'd378: r_data <= DATA_W'h00000000;
			DATA_W'd379: r_data <= DATA_W'h00000000;
			DATA_W'd380: r_data <= DATA_W'h00000000;
			DATA_W'd381: r_data <= DATA_W'h00000000;
			DATA_W'd382: r_data <= DATA_W'h00000000;
			DATA_W'd383: r_data <= DATA_W'h00000000;
			DATA_W'd384: r_data <= DATA_W'h00000000;
			DATA_W'd385: r_data <= DATA_W'h00000000;
			DATA_W'd386: r_data <= DATA_W'h00000000;
			DATA_W'd387: r_data <= DATA_W'h00000000;
			DATA_W'd388: r_data <= DATA_W'h00000000;
			DATA_W'd389: r_data <= DATA_W'h00000000;
			DATA_W'd390: r_data <= DATA_W'h00000000;
			DATA_W'd391: r_data <= DATA_W'h00000000;
			DATA_W'd392: r_data <= DATA_W'h00000000;
			DATA_W'd393: r_data <= DATA_W'h00000000;
			DATA_W'd394: r_data <= DATA_W'h00000000;
			DATA_W'd395: r_data <= DATA_W'h00000000;
			DATA_W'd396: r_data <= DATA_W'h00000000;
			DATA_W'd397: r_data <= DATA_W'h00000000;
			DATA_W'd398: r_data <= DATA_W'h00000000;
			DATA_W'd399: r_data <= DATA_W'h00000000;
			DATA_W'd400: r_data <= DATA_W'h00000000;
			DATA_W'd401: r_data <= DATA_W'h00000000;
			DATA_W'd402: r_data <= DATA_W'h00000000;
			DATA_W'd403: r_data <= DATA_W'h00000000;
			DATA_W'd404: r_data <= DATA_W'h00000000;
			DATA_W'd405: r_data <= DATA_W'h00000000;
			DATA_W'd406: r_data <= DATA_W'h00000000;
			DATA_W'd407: r_data <= DATA_W'h00000000;
			DATA_W'd408: r_data <= DATA_W'h00000000;
			DATA_W'd409: r_data <= DATA_W'h00000000;
			DATA_W'd410: r_data <= DATA_W'h00000000;
			DATA_W'd411: r_data <= DATA_W'h00000000;
			DATA_W'd412: r_data <= DATA_W'h00000000;
			DATA_W'd413: r_data <= DATA_W'h00000000;
			DATA_W'd414: r_data <= DATA_W'h00000000;
			DATA_W'd415: r_data <= DATA_W'h00000000;
			DATA_W'd416: r_data <= DATA_W'h00000000;
			DATA_W'd417: r_data <= DATA_W'h00000000;
			DATA_W'd418: r_data <= DATA_W'h00000000;
			DATA_W'd419: r_data <= DATA_W'h00000000;
			DATA_W'd420: r_data <= DATA_W'h00000000;
			DATA_W'd421: r_data <= DATA_W'h00000000;
			DATA_W'd422: r_data <= DATA_W'h00000000;
			DATA_W'd423: r_data <= DATA_W'h00000000;
			DATA_W'd424: r_data <= DATA_W'h00000000;
			DATA_W'd425: r_data <= DATA_W'h00000000;
			DATA_W'd426: r_data <= DATA_W'h00000000;
			DATA_W'd427: r_data <= DATA_W'h00000000;
			DATA_W'd428: r_data <= DATA_W'h00000000;
			DATA_W'd429: r_data <= DATA_W'h00000000;
			DATA_W'd430: r_data <= DATA_W'h00000000;
			DATA_W'd431: r_data <= DATA_W'h00000000;
			DATA_W'd432: r_data <= DATA_W'h00000000;
			DATA_W'd433: r_data <= DATA_W'h00000000;
			DATA_W'd434: r_data <= DATA_W'h00000000;
			DATA_W'd435: r_data <= DATA_W'h00000000;
			DATA_W'd436: r_data <= DATA_W'h00000000;
			DATA_W'd437: r_data <= DATA_W'h00000000;
			DATA_W'd438: r_data <= DATA_W'h00000000;
			DATA_W'd439: r_data <= DATA_W'h00000000;
			DATA_W'd440: r_data <= DATA_W'h00000000;
			DATA_W'd441: r_data <= DATA_W'h00000000;
			DATA_W'd442: r_data <= DATA_W'h00000000;
			DATA_W'd443: r_data <= DATA_W'h00000000;
			DATA_W'd444: r_data <= DATA_W'h00000000;
			DATA_W'd445: r_data <= DATA_W'h00000000;
			DATA_W'd446: r_data <= DATA_W'h00000000;
			DATA_W'd447: r_data <= DATA_W'h00000000;
			DATA_W'd448: r_data <= DATA_W'h00000000;
			DATA_W'd449: r_data <= DATA_W'h00000000;
			DATA_W'd450: r_data <= DATA_W'h00000000;
			DATA_W'd451: r_data <= DATA_W'h00000000;
			DATA_W'd452: r_data <= DATA_W'h00000000;
			DATA_W'd453: r_data <= DATA_W'h00000000;
			DATA_W'd454: r_data <= DATA_W'h00000000;
			DATA_W'd455: r_data <= DATA_W'h00000000;
			DATA_W'd456: r_data <= DATA_W'h00000000;
			DATA_W'd457: r_data <= DATA_W'h00000000;
			DATA_W'd458: r_data <= DATA_W'h00000000;
			DATA_W'd459: r_data <= DATA_W'h00000000;
			DATA_W'd460: r_data <= DATA_W'h00000000;
			DATA_W'd461: r_data <= DATA_W'h00000000;
			DATA_W'd462: r_data <= DATA_W'h00000000;
			DATA_W'd463: r_data <= DATA_W'h00000000;
			DATA_W'd464: r_data <= DATA_W'h00000000;
			DATA_W'd465: r_data <= DATA_W'h00000000;
			DATA_W'd466: r_data <= DATA_W'h00000000;
			DATA_W'd467: r_data <= DATA_W'h00000000;
			DATA_W'd468: r_data <= DATA_W'h00000000;
			DATA_W'd469: r_data <= DATA_W'h00000000;
			DATA_W'd470: r_data <= DATA_W'h00000000;
			DATA_W'd471: r_data <= DATA_W'h00000000;
			DATA_W'd472: r_data <= DATA_W'h00000000;
			DATA_W'd473: r_data <= DATA_W'h00000000;
			DATA_W'd474: r_data <= DATA_W'h00000000;
			DATA_W'd475: r_data <= DATA_W'h00000000;
			DATA_W'd476: r_data <= DATA_W'h00000000;
			DATA_W'd477: r_data <= DATA_W'h00000000;
			DATA_W'd478: r_data <= DATA_W'h00000000;
			DATA_W'd479: r_data <= DATA_W'h00000000;
			DATA_W'd480: r_data <= DATA_W'h00000000;
			DATA_W'd481: r_data <= DATA_W'h00000000;
			DATA_W'd482: r_data <= DATA_W'h00000000;
			DATA_W'd483: r_data <= DATA_W'h00000000;
			DATA_W'd484: r_data <= DATA_W'h00000000;
			DATA_W'd485: r_data <= DATA_W'h00000000;
			DATA_W'd486: r_data <= DATA_W'h00000000;
			DATA_W'd487: r_data <= DATA_W'h00000000;
			DATA_W'd488: r_data <= DATA_W'h00000000;
			DATA_W'd489: r_data <= DATA_W'h00000000;
			DATA_W'd490: r_data <= DATA_W'h00000000;
			DATA_W'd491: r_data <= DATA_W'h00000000;
			DATA_W'd492: r_data <= DATA_W'h00000000;
			DATA_W'd493: r_data <= DATA_W'h00000000;
			DATA_W'd494: r_data <= DATA_W'h00000000;
			DATA_W'd495: r_data <= DATA_W'h00000000;
			DATA_W'd496: r_data <= DATA_W'h00000000;
			DATA_W'd497: r_data <= DATA_W'h00000000;
			DATA_W'd498: r_data <= DATA_W'h00000000;
			DATA_W'd499: r_data <= DATA_W'h00000000;
			DATA_W'd500: r_data <= DATA_W'h00000000;
			DATA_W'd501: r_data <= DATA_W'h00000000;
			DATA_W'd502: r_data <= DATA_W'h00000000;
			DATA_W'd503: r_data <= DATA_W'h00000000;
			DATA_W'd504: r_data <= DATA_W'h00000000;
			DATA_W'd505: r_data <= DATA_W'h00000000;
			DATA_W'd506: r_data <= DATA_W'h00000000;
			DATA_W'd507: r_data <= DATA_W'h00000000;
			DATA_W'd508: r_data <= DATA_W'h00000000;
			DATA_W'd509: r_data <= DATA_W'h00000000;
			DATA_W'd510: r_data <= DATA_W'h00000000;
			DATA_W'd511: r_data <= DATA_W'h00000000;
			DATA_W'd512: r_data <= DATA_W'h00000000;
			DATA_W'd513: r_data <= DATA_W'h00000000;
			DATA_W'd514: r_data <= DATA_W'h00000000;
			DATA_W'd515: r_data <= DATA_W'h00000000;
			DATA_W'd516: r_data <= DATA_W'h00000000;
			DATA_W'd517: r_data <= DATA_W'h00000000;
			DATA_W'd518: r_data <= DATA_W'h00000000;
			DATA_W'd519: r_data <= DATA_W'h00000000;
			DATA_W'd520: r_data <= DATA_W'h00000000;
			DATA_W'd521: r_data <= DATA_W'h00000000;
			DATA_W'd522: r_data <= DATA_W'h00000000;
			DATA_W'd523: r_data <= DATA_W'h00000000;
			DATA_W'd524: r_data <= DATA_W'h00000000;
			DATA_W'd525: r_data <= DATA_W'h00000000;
			DATA_W'd526: r_data <= DATA_W'h00000000;
			DATA_W'd527: r_data <= DATA_W'h00000000;
			DATA_W'd528: r_data <= DATA_W'h00000000;
			DATA_W'd529: r_data <= DATA_W'h00000000;
			DATA_W'd530: r_data <= DATA_W'h00000000;
			DATA_W'd531: r_data <= DATA_W'h00000000;
			DATA_W'd532: r_data <= DATA_W'h00000000;
			DATA_W'd533: r_data <= DATA_W'h00000000;
			DATA_W'd534: r_data <= DATA_W'h00000000;
			DATA_W'd535: r_data <= DATA_W'h00000000;
			DATA_W'd536: r_data <= DATA_W'h00000000;
			DATA_W'd537: r_data <= DATA_W'h00000000;
			DATA_W'd538: r_data <= DATA_W'h00000000;
			DATA_W'd539: r_data <= DATA_W'h00000000;
			DATA_W'd540: r_data <= DATA_W'h00000000;
			DATA_W'd541: r_data <= DATA_W'h00000000;
			DATA_W'd542: r_data <= DATA_W'h00000000;
			DATA_W'd543: r_data <= DATA_W'h00000000;
			DATA_W'd544: r_data <= DATA_W'h00000000;
			DATA_W'd545: r_data <= DATA_W'h00000000;
			DATA_W'd546: r_data <= DATA_W'h00000000;
			DATA_W'd547: r_data <= DATA_W'h00000000;
			DATA_W'd548: r_data <= DATA_W'h00000000;
			DATA_W'd549: r_data <= DATA_W'h00000000;
			DATA_W'd550: r_data <= DATA_W'h00000000;
			DATA_W'd551: r_data <= DATA_W'h00000000;
			DATA_W'd552: r_data <= DATA_W'h00000000;
			DATA_W'd553: r_data <= DATA_W'h00000000;
			DATA_W'd554: r_data <= DATA_W'h00000000;
			DATA_W'd555: r_data <= DATA_W'h00000000;
			DATA_W'd556: r_data <= DATA_W'h00000000;
			DATA_W'd557: r_data <= DATA_W'h00000000;
			DATA_W'd558: r_data <= DATA_W'h00000000;
			DATA_W'd559: r_data <= DATA_W'h00000000;
			DATA_W'd560: r_data <= DATA_W'h00000000;
			DATA_W'd561: r_data <= DATA_W'h00000000;
			DATA_W'd562: r_data <= DATA_W'h00000000;
			DATA_W'd563: r_data <= DATA_W'h00000000;
			DATA_W'd564: r_data <= DATA_W'h00000000;
			DATA_W'd565: r_data <= DATA_W'h00000000;
			DATA_W'd566: r_data <= DATA_W'h00000000;
			DATA_W'd567: r_data <= DATA_W'h00000000;
			DATA_W'd568: r_data <= DATA_W'h00000000;
			DATA_W'd569: r_data <= DATA_W'h00000000;
			DATA_W'd570: r_data <= DATA_W'h00000000;
			DATA_W'd571: r_data <= DATA_W'h00000000;
			DATA_W'd572: r_data <= DATA_W'h00000000;
			DATA_W'd573: r_data <= DATA_W'h00000000;
			DATA_W'd574: r_data <= DATA_W'h00000000;
			DATA_W'd575: r_data <= DATA_W'h00000000;
			DATA_W'd576: r_data <= DATA_W'h00000000;
			DATA_W'd577: r_data <= DATA_W'h00000000;
			DATA_W'd578: r_data <= DATA_W'h00000000;
			DATA_W'd579: r_data <= DATA_W'h00000000;
			DATA_W'd580: r_data <= DATA_W'h00000000;
			DATA_W'd581: r_data <= DATA_W'h00000000;
			DATA_W'd582: r_data <= DATA_W'h00000000;
			DATA_W'd583: r_data <= DATA_W'h00000000;
			DATA_W'd584: r_data <= DATA_W'h00000000;
			DATA_W'd585: r_data <= DATA_W'h00000000;
			DATA_W'd586: r_data <= DATA_W'h00000000;
			DATA_W'd587: r_data <= DATA_W'h00000000;
			DATA_W'd588: r_data <= DATA_W'h00000000;
			DATA_W'd589: r_data <= DATA_W'h00000000;
			DATA_W'd590: r_data <= DATA_W'h00000000;
			DATA_W'd591: r_data <= DATA_W'h00000000;
			DATA_W'd592: r_data <= DATA_W'h00000000;
			DATA_W'd593: r_data <= DATA_W'h00000000;
			DATA_W'd594: r_data <= DATA_W'h00000000;
			DATA_W'd595: r_data <= DATA_W'h00000000;
			DATA_W'd596: r_data <= DATA_W'h00000000;
			DATA_W'd597: r_data <= DATA_W'h00000000;
			DATA_W'd598: r_data <= DATA_W'h00000000;
			DATA_W'd599: r_data <= DATA_W'h00000000;
			DATA_W'd600: r_data <= DATA_W'h00000000;
			DATA_W'd601: r_data <= DATA_W'h00000000;
			DATA_W'd602: r_data <= DATA_W'h00000000;
			DATA_W'd603: r_data <= DATA_W'h00000000;
			DATA_W'd604: r_data <= DATA_W'h00000000;
			DATA_W'd605: r_data <= DATA_W'h00000000;
			DATA_W'd606: r_data <= DATA_W'h00000000;
			DATA_W'd607: r_data <= DATA_W'h00000000;
			DATA_W'd608: r_data <= DATA_W'h00000000;
			DATA_W'd609: r_data <= DATA_W'h00000000;
			DATA_W'd610: r_data <= DATA_W'h00000000;
			DATA_W'd611: r_data <= DATA_W'h00000000;
			DATA_W'd612: r_data <= DATA_W'h00000000;
			DATA_W'd613: r_data <= DATA_W'h00000000;
			DATA_W'd614: r_data <= DATA_W'h00000000;
			DATA_W'd615: r_data <= DATA_W'h00000000;
			DATA_W'd616: r_data <= DATA_W'h00000000;
			DATA_W'd617: r_data <= DATA_W'h00000000;
			DATA_W'd618: r_data <= DATA_W'h00000000;
			DATA_W'd619: r_data <= DATA_W'h00000000;
			DATA_W'd620: r_data <= DATA_W'h00000000;
			DATA_W'd621: r_data <= DATA_W'h00000000;
			DATA_W'd622: r_data <= DATA_W'h00000000;
			DATA_W'd623: r_data <= DATA_W'h00000000;
			DATA_W'd624: r_data <= DATA_W'h00000000;
			DATA_W'd625: r_data <= DATA_W'h00000000;
			DATA_W'd626: r_data <= DATA_W'h00000000;
			DATA_W'd627: r_data <= DATA_W'h00000000;
			DATA_W'd628: r_data <= DATA_W'h00000000;
			DATA_W'd629: r_data <= DATA_W'h00000000;
			DATA_W'd630: r_data <= DATA_W'h00000000;
			DATA_W'd631: r_data <= DATA_W'h00000000;
			DATA_W'd632: r_data <= DATA_W'h00000000;
			DATA_W'd633: r_data <= DATA_W'h00000000;
			DATA_W'd634: r_data <= DATA_W'h00000000;
			DATA_W'd635: r_data <= DATA_W'h00000000;
			DATA_W'd636: r_data <= DATA_W'h00000000;
			DATA_W'd637: r_data <= DATA_W'h00000000;
			DATA_W'd638: r_data <= DATA_W'h00000000;
			DATA_W'd639: r_data <= DATA_W'h00000000;
			DATA_W'd640: r_data <= DATA_W'h00000000;
			DATA_W'd641: r_data <= DATA_W'h00000000;
			DATA_W'd642: r_data <= DATA_W'h00000000;
			DATA_W'd643: r_data <= DATA_W'h00000000;
			DATA_W'd644: r_data <= DATA_W'h00000000;
			DATA_W'd645: r_data <= DATA_W'h00000000;
			DATA_W'd646: r_data <= DATA_W'h00000000;
			DATA_W'd647: r_data <= DATA_W'h00000000;
			DATA_W'd648: r_data <= DATA_W'h00000000;
			DATA_W'd649: r_data <= DATA_W'h00000000;
			DATA_W'd650: r_data <= DATA_W'h00000000;
			DATA_W'd651: r_data <= DATA_W'h00000000;
			DATA_W'd652: r_data <= DATA_W'h00000000;
			DATA_W'd653: r_data <= DATA_W'h00000000;
			DATA_W'd654: r_data <= DATA_W'h00000000;
			DATA_W'd655: r_data <= DATA_W'h00000000;
			DATA_W'd656: r_data <= DATA_W'h00000000;
			DATA_W'd657: r_data <= DATA_W'h00000000;
			DATA_W'd658: r_data <= DATA_W'h00000000;
			DATA_W'd659: r_data <= DATA_W'h00000000;
			DATA_W'd660: r_data <= DATA_W'h00000000;
			DATA_W'd661: r_data <= DATA_W'h00000000;
			DATA_W'd662: r_data <= DATA_W'h00000000;
			DATA_W'd663: r_data <= DATA_W'h00000000;
			DATA_W'd664: r_data <= DATA_W'h00000000;
			DATA_W'd665: r_data <= DATA_W'h00000000;
			DATA_W'd666: r_data <= DATA_W'h00000000;
			DATA_W'd667: r_data <= DATA_W'h00000000;
			DATA_W'd668: r_data <= DATA_W'h00000000;
			DATA_W'd669: r_data <= DATA_W'h00000000;
			DATA_W'd670: r_data <= DATA_W'h00000000;
			DATA_W'd671: r_data <= DATA_W'h00000000;
			DATA_W'd672: r_data <= DATA_W'h00000000;
			DATA_W'd673: r_data <= DATA_W'h00000000;
			DATA_W'd674: r_data <= DATA_W'h00000000;
			DATA_W'd675: r_data <= DATA_W'h00000000;
			DATA_W'd676: r_data <= DATA_W'h00000000;
			DATA_W'd677: r_data <= DATA_W'h00000000;
			DATA_W'd678: r_data <= DATA_W'h00000000;
			DATA_W'd679: r_data <= DATA_W'h00000000;
			DATA_W'd680: r_data <= DATA_W'h00000000;
			DATA_W'd681: r_data <= DATA_W'h00000000;
			DATA_W'd682: r_data <= DATA_W'h00000000;
			DATA_W'd683: r_data <= DATA_W'h00000000;
			DATA_W'd684: r_data <= DATA_W'h00000000;
			DATA_W'd685: r_data <= DATA_W'h00000000;
			DATA_W'd686: r_data <= DATA_W'h00000000;
			DATA_W'd687: r_data <= DATA_W'h00000000;
			DATA_W'd688: r_data <= DATA_W'h00000000;
			DATA_W'd689: r_data <= DATA_W'h00000000;
			DATA_W'd690: r_data <= DATA_W'h00000000;
			DATA_W'd691: r_data <= DATA_W'h00000000;
			DATA_W'd692: r_data <= DATA_W'h00000000;
			DATA_W'd693: r_data <= DATA_W'h00000000;
			DATA_W'd694: r_data <= DATA_W'h00000000;
			DATA_W'd695: r_data <= DATA_W'h00000000;
			DATA_W'd696: r_data <= DATA_W'h00000000;
			DATA_W'd697: r_data <= DATA_W'h00000000;
			DATA_W'd698: r_data <= DATA_W'h00000000;
			DATA_W'd699: r_data <= DATA_W'h00000000;
			DATA_W'd700: r_data <= DATA_W'h00000000;
			DATA_W'd701: r_data <= DATA_W'h00000000;
			DATA_W'd702: r_data <= DATA_W'h00000000;
			DATA_W'd703: r_data <= DATA_W'h00000000;
			DATA_W'd704: r_data <= DATA_W'h00000000;
			DATA_W'd705: r_data <= DATA_W'h00000000;
			DATA_W'd706: r_data <= DATA_W'h00000000;
			DATA_W'd707: r_data <= DATA_W'h00000000;
			DATA_W'd708: r_data <= DATA_W'h00000000;
			DATA_W'd709: r_data <= DATA_W'h00000000;
			DATA_W'd710: r_data <= DATA_W'h00000000;
			DATA_W'd711: r_data <= DATA_W'h00000000;
			DATA_W'd712: r_data <= DATA_W'h00000000;
			DATA_W'd713: r_data <= DATA_W'h00000000;
			DATA_W'd714: r_data <= DATA_W'h00000000;
			DATA_W'd715: r_data <= DATA_W'h00000000;
			DATA_W'd716: r_data <= DATA_W'h00000000;
			DATA_W'd717: r_data <= DATA_W'h00000000;
			DATA_W'd718: r_data <= DATA_W'h00000000;
			DATA_W'd719: r_data <= DATA_W'h00000000;
			DATA_W'd720: r_data <= DATA_W'h00000000;
			DATA_W'd721: r_data <= DATA_W'h00000000;
			DATA_W'd722: r_data <= DATA_W'h00000000;
			DATA_W'd723: r_data <= DATA_W'h00000000;
			DATA_W'd724: r_data <= DATA_W'h00000000;
			DATA_W'd725: r_data <= DATA_W'h00000000;
			DATA_W'd726: r_data <= DATA_W'h00000000;
			DATA_W'd727: r_data <= DATA_W'h00000000;
			DATA_W'd728: r_data <= DATA_W'h00000000;
			DATA_W'd729: r_data <= DATA_W'h00000000;
			DATA_W'd730: r_data <= DATA_W'h00000000;
			DATA_W'd731: r_data <= DATA_W'h00000000;
			DATA_W'd732: r_data <= DATA_W'h00000000;
			DATA_W'd733: r_data <= DATA_W'h00000000;
			DATA_W'd734: r_data <= DATA_W'h00000000;
			DATA_W'd735: r_data <= DATA_W'h00000000;
			DATA_W'd736: r_data <= DATA_W'h00000000;
			DATA_W'd737: r_data <= DATA_W'h00000000;
			DATA_W'd738: r_data <= DATA_W'h00000000;
			DATA_W'd739: r_data <= DATA_W'h00000000;
			DATA_W'd740: r_data <= DATA_W'h00000000;
			DATA_W'd741: r_data <= DATA_W'h00000000;
			DATA_W'd742: r_data <= DATA_W'h00000000;
			DATA_W'd743: r_data <= DATA_W'h00000000;
			DATA_W'd744: r_data <= DATA_W'h00000000;
			DATA_W'd745: r_data <= DATA_W'h00000000;
			DATA_W'd746: r_data <= DATA_W'h00000000;
			DATA_W'd747: r_data <= DATA_W'h00000000;
			DATA_W'd748: r_data <= DATA_W'h00000000;
			DATA_W'd749: r_data <= DATA_W'h00000000;
			DATA_W'd750: r_data <= DATA_W'h00000000;
			DATA_W'd751: r_data <= DATA_W'h00000000;
			DATA_W'd752: r_data <= DATA_W'h00000000;
			DATA_W'd753: r_data <= DATA_W'h00000000;
			DATA_W'd754: r_data <= DATA_W'h00000000;
			DATA_W'd755: r_data <= DATA_W'h00000000;
			DATA_W'd756: r_data <= DATA_W'h00000000;
			DATA_W'd757: r_data <= DATA_W'h00000000;
			DATA_W'd758: r_data <= DATA_W'h00000000;
			DATA_W'd759: r_data <= DATA_W'h00000000;
			DATA_W'd760: r_data <= DATA_W'h00000000;
			DATA_W'd761: r_data <= DATA_W'h00000000;
			DATA_W'd762: r_data <= DATA_W'h00000000;
			DATA_W'd763: r_data <= DATA_W'h00000000;
			DATA_W'd764: r_data <= DATA_W'h00000000;
			DATA_W'd765: r_data <= DATA_W'h00000000;
			DATA_W'd766: r_data <= DATA_W'h00000000;
			DATA_W'd767: r_data <= DATA_W'h00000000;
			DATA_W'd768: r_data <= DATA_W'h00000000;
			DATA_W'd769: r_data <= DATA_W'h00000000;
			DATA_W'd770: r_data <= DATA_W'h00000000;
			DATA_W'd771: r_data <= DATA_W'h00000000;
			DATA_W'd772: r_data <= DATA_W'h00000000;
			DATA_W'd773: r_data <= DATA_W'h00000000;
			DATA_W'd774: r_data <= DATA_W'h00000000;
			DATA_W'd775: r_data <= DATA_W'h00000000;
			DATA_W'd776: r_data <= DATA_W'h00000000;
			DATA_W'd777: r_data <= DATA_W'h00000000;
			DATA_W'd778: r_data <= DATA_W'h00000000;
			DATA_W'd779: r_data <= DATA_W'h00000000;
			DATA_W'd780: r_data <= DATA_W'h00000000;
			DATA_W'd781: r_data <= DATA_W'h00000000;
			DATA_W'd782: r_data <= DATA_W'h00000000;
			DATA_W'd783: r_data <= DATA_W'h00000000;
			DATA_W'd784: r_data <= DATA_W'h00000000;
			DATA_W'd785: r_data <= DATA_W'h00000000;
			DATA_W'd786: r_data <= DATA_W'h00000000;
			DATA_W'd787: r_data <= DATA_W'h00000000;
			DATA_W'd788: r_data <= DATA_W'h00000000;
			DATA_W'd789: r_data <= DATA_W'h00000000;
			DATA_W'd790: r_data <= DATA_W'h00000000;
			DATA_W'd791: r_data <= DATA_W'h00000000;
			DATA_W'd792: r_data <= DATA_W'h00000000;
			DATA_W'd793: r_data <= DATA_W'h00000000;
			DATA_W'd794: r_data <= DATA_W'h00000000;
			DATA_W'd795: r_data <= DATA_W'h00000000;
			DATA_W'd796: r_data <= DATA_W'h00000000;
			DATA_W'd797: r_data <= DATA_W'h00000000;
			DATA_W'd798: r_data <= DATA_W'h00000000;
			DATA_W'd799: r_data <= DATA_W'h00000000;
			DATA_W'd800: r_data <= DATA_W'h00000000;
			DATA_W'd801: r_data <= DATA_W'h00000000;
			DATA_W'd802: r_data <= DATA_W'h00000000;
			DATA_W'd803: r_data <= DATA_W'h00000000;
			DATA_W'd804: r_data <= DATA_W'h00000000;
			DATA_W'd805: r_data <= DATA_W'h00000000;
			DATA_W'd806: r_data <= DATA_W'h00000000;
			DATA_W'd807: r_data <= DATA_W'h00000000;
			DATA_W'd808: r_data <= DATA_W'h00000000;
			DATA_W'd809: r_data <= DATA_W'h00000000;
			DATA_W'd810: r_data <= DATA_W'h00000000;
			DATA_W'd811: r_data <= DATA_W'h00000000;
			DATA_W'd812: r_data <= DATA_W'h00000000;
			DATA_W'd813: r_data <= DATA_W'h00000000;
			DATA_W'd814: r_data <= DATA_W'h00000000;
			DATA_W'd815: r_data <= DATA_W'h00000000;
			DATA_W'd816: r_data <= DATA_W'h00000000;
			DATA_W'd817: r_data <= DATA_W'h00000000;
			DATA_W'd818: r_data <= DATA_W'h00000000;
			DATA_W'd819: r_data <= DATA_W'h00000000;
			DATA_W'd820: r_data <= DATA_W'h00000000;
			DATA_W'd821: r_data <= DATA_W'h00000000;
			DATA_W'd822: r_data <= DATA_W'h00000000;
			DATA_W'd823: r_data <= DATA_W'h00000000;
			DATA_W'd824: r_data <= DATA_W'h00000000;
			DATA_W'd825: r_data <= DATA_W'h00000000;
			DATA_W'd826: r_data <= DATA_W'h00000000;
			DATA_W'd827: r_data <= DATA_W'h00000000;
			DATA_W'd828: r_data <= DATA_W'h00000000;
			DATA_W'd829: r_data <= DATA_W'h00000000;
			DATA_W'd830: r_data <= DATA_W'h00000000;
			DATA_W'd831: r_data <= DATA_W'h00000000;
			DATA_W'd832: r_data <= DATA_W'h00000000;
			DATA_W'd833: r_data <= DATA_W'h00000000;
			DATA_W'd834: r_data <= DATA_W'h00000000;
			DATA_W'd835: r_data <= DATA_W'h00000000;
			DATA_W'd836: r_data <= DATA_W'h00000000;
			DATA_W'd837: r_data <= DATA_W'h00000000;
			DATA_W'd838: r_data <= DATA_W'h00000000;
			DATA_W'd839: r_data <= DATA_W'h00000000;
			DATA_W'd840: r_data <= DATA_W'h00000000;
			DATA_W'd841: r_data <= DATA_W'h00000000;
			DATA_W'd842: r_data <= DATA_W'h00000000;
			DATA_W'd843: r_data <= DATA_W'h00000000;
			DATA_W'd844: r_data <= DATA_W'h00000000;
			DATA_W'd845: r_data <= DATA_W'h00000000;
			DATA_W'd846: r_data <= DATA_W'h00000000;
			DATA_W'd847: r_data <= DATA_W'h00000000;
			DATA_W'd848: r_data <= DATA_W'h00000000;
			DATA_W'd849: r_data <= DATA_W'h00000000;
			DATA_W'd850: r_data <= DATA_W'h00000000;
			DATA_W'd851: r_data <= DATA_W'h00000000;
			DATA_W'd852: r_data <= DATA_W'h00000000;
			DATA_W'd853: r_data <= DATA_W'h00000000;
			DATA_W'd854: r_data <= DATA_W'h00000000;
			DATA_W'd855: r_data <= DATA_W'h00000000;
			DATA_W'd856: r_data <= DATA_W'h00000000;
			DATA_W'd857: r_data <= DATA_W'h00000000;
			DATA_W'd858: r_data <= DATA_W'h00000000;
			DATA_W'd859: r_data <= DATA_W'h00000000;
			DATA_W'd860: r_data <= DATA_W'h00000000;
			DATA_W'd861: r_data <= DATA_W'h00000000;
			DATA_W'd862: r_data <= DATA_W'h00000000;
			DATA_W'd863: r_data <= DATA_W'h00000000;
			DATA_W'd864: r_data <= DATA_W'h00000000;
			DATA_W'd865: r_data <= DATA_W'h00000000;
			DATA_W'd866: r_data <= DATA_W'h00000000;
			DATA_W'd867: r_data <= DATA_W'h00000000;
			DATA_W'd868: r_data <= DATA_W'h00000000;
			DATA_W'd869: r_data <= DATA_W'h00000000;
			DATA_W'd870: r_data <= DATA_W'h00000000;
			DATA_W'd871: r_data <= DATA_W'h00000000;
			DATA_W'd872: r_data <= DATA_W'h00000000;
			DATA_W'd873: r_data <= DATA_W'h00000000;
			DATA_W'd874: r_data <= DATA_W'h00000000;
			DATA_W'd875: r_data <= DATA_W'h00000000;
			DATA_W'd876: r_data <= DATA_W'h00000000;
			DATA_W'd877: r_data <= DATA_W'h00000000;
			DATA_W'd878: r_data <= DATA_W'h00000000;
			DATA_W'd879: r_data <= DATA_W'h00000000;
			DATA_W'd880: r_data <= DATA_W'h00000000;
			DATA_W'd881: r_data <= DATA_W'h00000000;
			DATA_W'd882: r_data <= DATA_W'h00000000;
			DATA_W'd883: r_data <= DATA_W'h00000000;
			DATA_W'd884: r_data <= DATA_W'h00000000;
			DATA_W'd885: r_data <= DATA_W'h00000000;
			DATA_W'd886: r_data <= DATA_W'h00000000;
			DATA_W'd887: r_data <= DATA_W'h00000000;
			DATA_W'd888: r_data <= DATA_W'h00000000;
			DATA_W'd889: r_data <= DATA_W'h00000000;
			DATA_W'd890: r_data <= DATA_W'h00000000;
			DATA_W'd891: r_data <= DATA_W'h00000000;
			DATA_W'd892: r_data <= DATA_W'h00000000;
			DATA_W'd893: r_data <= DATA_W'h00000000;
			DATA_W'd894: r_data <= DATA_W'h00000000;
			DATA_W'd895: r_data <= DATA_W'h00000000;
			DATA_W'd896: r_data <= DATA_W'h00000000;
			DATA_W'd897: r_data <= DATA_W'h00000000;
			DATA_W'd898: r_data <= DATA_W'h00000000;
			DATA_W'd899: r_data <= DATA_W'h00000000;
			DATA_W'd900: r_data <= DATA_W'h00000000;
			DATA_W'd901: r_data <= DATA_W'h00000000;
			DATA_W'd902: r_data <= DATA_W'h00000000;
			DATA_W'd903: r_data <= DATA_W'h00000000;
			DATA_W'd904: r_data <= DATA_W'h00000000;
			DATA_W'd905: r_data <= DATA_W'h00000000;
			DATA_W'd906: r_data <= DATA_W'h00000000;
			DATA_W'd907: r_data <= DATA_W'h00000000;
			DATA_W'd908: r_data <= DATA_W'h00000000;
			DATA_W'd909: r_data <= DATA_W'h00000000;
			DATA_W'd910: r_data <= DATA_W'h00000000;
			DATA_W'd911: r_data <= DATA_W'h00000000;
			DATA_W'd912: r_data <= DATA_W'h00000000;
			DATA_W'd913: r_data <= DATA_W'h00000000;
			DATA_W'd914: r_data <= DATA_W'h00000000;
			DATA_W'd915: r_data <= DATA_W'h00000000;
			DATA_W'd916: r_data <= DATA_W'h00000000;
			DATA_W'd917: r_data <= DATA_W'h00000000;
			DATA_W'd918: r_data <= DATA_W'h00000000;
			DATA_W'd919: r_data <= DATA_W'h00000000;
			DATA_W'd920: r_data <= DATA_W'h00000000;
			DATA_W'd921: r_data <= DATA_W'h00000000;
			DATA_W'd922: r_data <= DATA_W'h00000000;
			DATA_W'd923: r_data <= DATA_W'h00000000;
			DATA_W'd924: r_data <= DATA_W'h00000000;
			DATA_W'd925: r_data <= DATA_W'h00000000;
			DATA_W'd926: r_data <= DATA_W'h00000000;
			DATA_W'd927: r_data <= DATA_W'h00000000;
			DATA_W'd928: r_data <= DATA_W'h00000000;
			DATA_W'd929: r_data <= DATA_W'h00000000;
			DATA_W'd930: r_data <= DATA_W'h00000000;
			DATA_W'd931: r_data <= DATA_W'h00000000;
			DATA_W'd932: r_data <= DATA_W'h00000000;
			DATA_W'd933: r_data <= DATA_W'h00000000;
			DATA_W'd934: r_data <= DATA_W'h00000000;
			DATA_W'd935: r_data <= DATA_W'h00000000;
			DATA_W'd936: r_data <= DATA_W'h00000000;
			DATA_W'd937: r_data <= DATA_W'h00000000;
			DATA_W'd938: r_data <= DATA_W'h00000000;
			DATA_W'd939: r_data <= DATA_W'h00000000;
			DATA_W'd940: r_data <= DATA_W'h00000000;
			DATA_W'd941: r_data <= DATA_W'h00000000;
			DATA_W'd942: r_data <= DATA_W'h00000000;
			DATA_W'd943: r_data <= DATA_W'h00000000;
			DATA_W'd944: r_data <= DATA_W'h00000000;
			DATA_W'd945: r_data <= DATA_W'h00000000;
			DATA_W'd946: r_data <= DATA_W'h00000000;
			DATA_W'd947: r_data <= DATA_W'h00000000;
			DATA_W'd948: r_data <= DATA_W'h00000000;
			DATA_W'd949: r_data <= DATA_W'h00000000;
			DATA_W'd950: r_data <= DATA_W'h00000000;
			DATA_W'd951: r_data <= DATA_W'h00000000;
			DATA_W'd952: r_data <= DATA_W'h00000000;
			DATA_W'd953: r_data <= DATA_W'h00000000;
			DATA_W'd954: r_data <= DATA_W'h00000000;
			DATA_W'd955: r_data <= DATA_W'h00000000;
			DATA_W'd956: r_data <= DATA_W'h00000000;
			DATA_W'd957: r_data <= DATA_W'h00000000;
			DATA_W'd958: r_data <= DATA_W'h00000000;
			DATA_W'd959: r_data <= DATA_W'h00000000;
			DATA_W'd960: r_data <= DATA_W'h00000000;
			DATA_W'd961: r_data <= DATA_W'h00000000;
			DATA_W'd962: r_data <= DATA_W'h00000000;
			DATA_W'd963: r_data <= DATA_W'h00000000;
			DATA_W'd964: r_data <= DATA_W'h00000000;
			DATA_W'd965: r_data <= DATA_W'h00000000;
			DATA_W'd966: r_data <= DATA_W'h00000000;
			DATA_W'd967: r_data <= DATA_W'h00000000;
			DATA_W'd968: r_data <= DATA_W'h00000000;
			DATA_W'd969: r_data <= DATA_W'h00000000;
			DATA_W'd970: r_data <= DATA_W'h00000000;
			DATA_W'd971: r_data <= DATA_W'h00000000;
			DATA_W'd972: r_data <= DATA_W'h00000000;
			DATA_W'd973: r_data <= DATA_W'h00000000;
			DATA_W'd974: r_data <= DATA_W'h00000000;
			DATA_W'd975: r_data <= DATA_W'h00000000;
			DATA_W'd976: r_data <= DATA_W'h00000000;
			DATA_W'd977: r_data <= DATA_W'h00000000;
			DATA_W'd978: r_data <= DATA_W'h00000000;
			DATA_W'd979: r_data <= DATA_W'h00000000;
			DATA_W'd980: r_data <= DATA_W'h00000000;
			DATA_W'd981: r_data <= DATA_W'h00000000;
			DATA_W'd982: r_data <= DATA_W'h00000000;
			DATA_W'd983: r_data <= DATA_W'h00000000;
			DATA_W'd984: r_data <= DATA_W'h00000000;
			DATA_W'd985: r_data <= DATA_W'h00000000;
			DATA_W'd986: r_data <= DATA_W'h00000000;
			DATA_W'd987: r_data <= DATA_W'h00000000;
			DATA_W'd988: r_data <= DATA_W'h00000000;
			DATA_W'd989: r_data <= DATA_W'h00000000;
			DATA_W'd990: r_data <= DATA_W'h00000000;
			DATA_W'd991: r_data <= DATA_W'h00000000;
			DATA_W'd992: r_data <= DATA_W'h00000000;
			DATA_W'd993: r_data <= DATA_W'h00000000;
			DATA_W'd994: r_data <= DATA_W'h00000000;
			DATA_W'd995: r_data <= DATA_W'h00000000;
			DATA_W'd996: r_data <= DATA_W'h00000000;
			DATA_W'd997: r_data <= DATA_W'h00000000;
			DATA_W'd998: r_data <= DATA_W'h00000000;
			DATA_W'd999: r_data <= DATA_W'h00000000;
			DATA_W'd1000: r_data <= DATA_W'h00000000;
			DATA_W'd1001: r_data <= DATA_W'h00000000;
			DATA_W'd1002: r_data <= DATA_W'h00000000;
			DATA_W'd1003: r_data <= DATA_W'h00000000;
			DATA_W'd1004: r_data <= DATA_W'h00000000;
			DATA_W'd1005: r_data <= DATA_W'h00000000;
			DATA_W'd1006: r_data <= DATA_W'h00000000;
			DATA_W'd1007: r_data <= DATA_W'h00000000;
			DATA_W'd1008: r_data <= DATA_W'h00000000;
			DATA_W'd1009: r_data <= DATA_W'h00000000;
			DATA_W'd1010: r_data <= DATA_W'h00000000;
			DATA_W'd1011: r_data <= DATA_W'h00000000;
			DATA_W'd1012: r_data <= DATA_W'h00000000;
			DATA_W'd1013: r_data <= DATA_W'h00000000;
			DATA_W'd1014: r_data <= DATA_W'h00000000;
			DATA_W'd1015: r_data <= DATA_W'h00000000;
			DATA_W'd1016: r_data <= DATA_W'h00000000;
			DATA_W'd1017: r_data <= DATA_W'h00000000;
			DATA_W'd1018: r_data <= DATA_W'h00000000;
			DATA_W'd1019: r_data <= DATA_W'h00000000;
			DATA_W'd1020: r_data <= DATA_W'h00000000;
			DATA_W'd1021: r_data <= DATA_W'h00000000;
			DATA_W'd1022: r_data <= DATA_W'h00000000;
			DATA_W'd1023: r_data <= DATA_W'h00000000;
			default: r_data <= DATA_W'h0;
		endcase
	end
